`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/21/2025 11:05:37 AM
// Design Name: 
// Module Name: matrix_mul64x10
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module multi_7x41( // 41 bit and 7 bti
input logic clk,rst,
input logic signed  [47:0] mul2_A, 
input logic signed [8:0] mul2_B,
output logic signed [55:0] mul2_res // 49 bit without sign
);
assign mul2_res = mul2_A*mul2_B;
endmodule


module adder_64in(
input logic clk,rst,
input logic signed [55:0] in_A1_0,  
 input logic signed [55:0] in_A1_1,   
 input logic signed [55:0] in_A1_2,   
 input logic signed [55:0] in_A1_3,   
 input logic signed [55:0] in_A1_4,   
 input logic signed [55:0] in_A1_5,   
 input logic signed [55:0] in_A1_6,   
 input logic signed [55:0] in_A1_7,   
 input logic signed [55:0] in_A1_8,   
 input logic signed [55:0] in_A1_9,   
 input logic signed [55:0] in_A1_10,  
 input logic signed [55:0] in_A1_11,  
 input logic signed [55:0] in_A1_12,  
 input logic signed [55:0] in_A1_13,  
 input logic signed [55:0] in_A1_14,  
 input logic signed [55:0] in_A1_15,  
 input logic signed [55:0] in_A1_16,  
 input logic signed [55:0] in_A1_17,  
 input logic signed [55:0] in_A1_18,
 input logic signed [55:0] in_A1_19,
 input logic signed [55:0] in_A1_20,
 input logic signed [55:0] in_A1_21,
 input logic signed [55:0] in_A1_22,
 input logic signed [55:0] in_A1_23,
 input logic signed [55:0] in_A1_24,
 input logic signed [55:0] in_A1_25,
 input logic signed [55:0] in_A1_26,
 input logic signed [55:0] in_A1_27,
 input logic signed [55:0] in_A1_28,
 input logic signed [55:0] in_A1_29,
 input logic signed [55:0] in_A1_30,
 input logic signed [55:0] in_A1_31,
 input logic signed [55:0] in_A1_32,
 input logic signed [55:0] in_A1_33,
 input logic signed [55:0] in_A1_34,
 input logic signed [55:0] in_A1_35,
 input logic signed [55:0] in_A1_36,
 input logic signed [55:0] in_A1_37,
 input logic signed [55:0] in_A1_38,
 input logic signed [55:0] in_A1_39,
 input logic signed [55:0] in_A1_40,
 input logic signed [55:0] in_A1_41,
 input logic signed [55:0] in_A1_42,
 input logic signed [55:0] in_A1_43,
 input logic signed [55:0] in_A1_44,
 input logic signed [55:0] in_A1_45,
 input logic signed [55:0] in_A1_46,
 input logic signed [55:0] in_A1_47,
 input logic signed [55:0] in_A1_48,
 input logic signed [55:0] in_A1_49,
 input logic signed [55:0] in_A1_50,
 input logic signed [55:0] in_A1_51,
 input logic signed [55:0] in_A1_52,
 input logic signed [55:0] in_A1_53,
 input logic signed [55:0] in_A1_54,
 input logic signed [55:0] in_A1_55,
 input logic signed [55:0] in_A1_56,
 input logic signed [55:0] in_A1_57,
 input logic signed [55:0] in_A1_58,
 input logic signed [55:0] in_A1_59,
 input logic signed [55:0] in_A1_60,
 input logic signed [55:0] in_A1_61,
 input logic signed [55:0] in_A1_62,
 input logic signed [55:0] in_A1_63,
output logic signed [61:0] out2_A 
    );
    
    assign  out2_A = in_A1_0 +  in_A1_1 +  in_A1_2 +  in_A1_3 +  in_A1_4 +  in_A1_5 +  in_A1_6 +  in_A1_7 +  in_A1_8 +  in_A1_9 +  in_A1_10 +  in_A1_11 +  in_A1_12 +  in_A1_13 +  in_A1_14 +  in_A1_15 +  in_A1_16 +  in_A1_17
     +  in_A1_18 +  in_A1_19 +  in_A1_20 +  in_A1_21 +  in_A1_22 +  in_A1_23 +  in_A1_24 +  in_A1_25 +  in_A1_26 +  in_A1_27 +  in_A1_28 +  in_A1_29 +  in_A1_30 +  in_A1_31 +  in_A1_32 +  in_A1_33 +  in_A1_34 +  in_A1_35 
     +  in_A1_36 +  in_A1_37 +  in_A1_38 +  in_A1_39 +  in_A1_40 +  in_A1_41 +  in_A1_42 +  in_A1_43 +  in_A1_44 +  in_A1_45 +  in_A1_46 +  in_A1_47 +  in_A1_48 +  in_A1_49 +  in_A1_50 +  in_A1_51 +  in_A1_52 +  in_A1_53 
     +  in_A1_54 +  in_A1_55 +  in_A1_56 +  in_A1_57 +  in_A1_58 +  in_A1_59 +  in_A1_60 +  in_A1_61 +  in_A1_62 +  in_A1_63;
endmodule



module matrix_mul64x10 (
input logic clk,rst,
input logic signed [47:0]matrix2_A [0:63], // flattened  
input logic signed [8:0]matrix2_B [0:639], //10*64
output logic signed[61:0] result_fc2 [0:9]
);


logic [55:0] mul_res2 [0:639];



multi_7x41 multi_7x41_mod_0(clk,rst,matrix2_A[0],matrix2_B[0],mul_res2[0]);
multi_7x41 multi_7x41_mod_1(clk,rst,matrix2_A[1],matrix2_B[1],mul_res2[1]);    
multi_7x41 multi_7x41_mod_2(clk,rst,matrix2_A[2],matrix2_B[2],mul_res2[2]);    
multi_7x41 multi_7x41_mod_3(clk,rst,matrix2_A[3],matrix2_B[3],mul_res2[3]);    
multi_7x41 multi_7x41_mod_4(clk,rst,matrix2_A[4],matrix2_B[4],mul_res2[4]);    
multi_7x41 multi_7x41_mod_5(clk,rst,matrix2_A[5],matrix2_B[5],mul_res2[5]);    
multi_7x41 multi_7x41_mod_6(clk,rst,matrix2_A[6],matrix2_B[6],mul_res2[6]);    
multi_7x41 multi_7x41_mod_7(clk,rst,matrix2_A[7],matrix2_B[7],mul_res2[7]);    
multi_7x41 multi_7x41_mod_8(clk,rst,matrix2_A[8],matrix2_B[8],mul_res2[8]);    
multi_7x41 multi_7x41_mod_9(clk,rst,matrix2_A[9],matrix2_B[9],mul_res2[9]);    
multi_7x41 multi_7x41_mod_10(clk,rst,matrix2_A[10],matrix2_B[10],mul_res2[10]);
multi_7x41 multi_7x41_mod_11(clk,rst,matrix2_A[11],matrix2_B[11],mul_res2[11]);
multi_7x41 multi_7x41_mod_12(clk,rst,matrix2_A[12],matrix2_B[12],mul_res2[12]);
multi_7x41 multi_7x41_mod_13(clk,rst,matrix2_A[13],matrix2_B[13],mul_res2[13]);
multi_7x41 multi_7x41_mod_14(clk,rst,matrix2_A[14],matrix2_B[14],mul_res2[14]);
multi_7x41 multi_7x41_mod_15(clk,rst,matrix2_A[15],matrix2_B[15],mul_res2[15]);
multi_7x41 multi_7x41_mod_16(clk,rst,matrix2_A[16],matrix2_B[16],mul_res2[16]);
multi_7x41 multi_7x41_mod_17(clk,rst,matrix2_A[17],matrix2_B[17],mul_res2[17]);
multi_7x41 multi_7x41_mod_18(clk,rst,matrix2_A[18],matrix2_B[18],mul_res2[18]);
multi_7x41 multi_7x41_mod_19(clk,rst,matrix2_A[19],matrix2_B[19],mul_res2[19]);
multi_7x41 multi_7x41_mod_20(clk,rst,matrix2_A[20],matrix2_B[20],mul_res2[20]);
multi_7x41 multi_7x41_mod_21(clk,rst,matrix2_A[21],matrix2_B[21],mul_res2[21]);
multi_7x41 multi_7x41_mod_22(clk,rst,matrix2_A[22],matrix2_B[22],mul_res2[22]);
multi_7x41 multi_7x41_mod_23(clk,rst,matrix2_A[23],matrix2_B[23],mul_res2[23]);
multi_7x41 multi_7x41_mod_24(clk,rst,matrix2_A[24],matrix2_B[24],mul_res2[24]);
multi_7x41 multi_7x41_mod_25(clk,rst,matrix2_A[25],matrix2_B[25],mul_res2[25]);
multi_7x41 multi_7x41_mod_26(clk,rst,matrix2_A[26],matrix2_B[26],mul_res2[26]);
multi_7x41 multi_7x41_mod_27(clk,rst,matrix2_A[27],matrix2_B[27],mul_res2[27]);
multi_7x41 multi_7x41_mod_28(clk,rst,matrix2_A[28],matrix2_B[28],mul_res2[28]);
multi_7x41 multi_7x41_mod_29(clk,rst,matrix2_A[29],matrix2_B[29],mul_res2[29]);
multi_7x41 multi_7x41_mod_30(clk,rst,matrix2_A[30],matrix2_B[30],mul_res2[30]);
multi_7x41 multi_7x41_mod_31(clk,rst,matrix2_A[31],matrix2_B[31],mul_res2[31]);
multi_7x41 multi_7x41_mod_32(clk,rst,matrix2_A[32],matrix2_B[32],mul_res2[32]);
multi_7x41 multi_7x41_mod_33(clk,rst,matrix2_A[33],matrix2_B[33],mul_res2[33]);
multi_7x41 multi_7x41_mod_34(clk,rst,matrix2_A[34],matrix2_B[34],mul_res2[34]);
multi_7x41 multi_7x41_mod_35(clk,rst,matrix2_A[35],matrix2_B[35],mul_res2[35]);
multi_7x41 multi_7x41_mod_36(clk,rst,matrix2_A[36],matrix2_B[36],mul_res2[36]);
multi_7x41 multi_7x41_mod_37(clk,rst,matrix2_A[37],matrix2_B[37],mul_res2[37]);
multi_7x41 multi_7x41_mod_38(clk,rst,matrix2_A[38],matrix2_B[38],mul_res2[38]);
multi_7x41 multi_7x41_mod_39(clk,rst,matrix2_A[39],matrix2_B[39],mul_res2[39]);
multi_7x41 multi_7x41_mod_40(clk,rst,matrix2_A[40],matrix2_B[40],mul_res2[40]);
multi_7x41 multi_7x41_mod_41(clk,rst,matrix2_A[41],matrix2_B[41],mul_res2[41]);
multi_7x41 multi_7x41_mod_42(clk,rst,matrix2_A[42],matrix2_B[42],mul_res2[42]);
multi_7x41 multi_7x41_mod_43(clk,rst,matrix2_A[43],matrix2_B[43],mul_res2[43]);
multi_7x41 multi_7x41_mod_44(clk,rst,matrix2_A[44],matrix2_B[44],mul_res2[44]);
multi_7x41 multi_7x41_mod_45(clk,rst,matrix2_A[45],matrix2_B[45],mul_res2[45]);
multi_7x41 multi_7x41_mod_46(clk,rst,matrix2_A[46],matrix2_B[46],mul_res2[46]);
multi_7x41 multi_7x41_mod_47(clk,rst,matrix2_A[47],matrix2_B[47],mul_res2[47]);
multi_7x41 multi_7x41_mod_48(clk,rst,matrix2_A[48],matrix2_B[48],mul_res2[48]);
multi_7x41 multi_7x41_mod_49(clk,rst,matrix2_A[49],matrix2_B[49],mul_res2[49]);
multi_7x41 multi_7x41_mod_50(clk,rst,matrix2_A[50],matrix2_B[50],mul_res2[50]);
multi_7x41 multi_7x41_mod_51(clk,rst,matrix2_A[51],matrix2_B[51],mul_res2[51]);
multi_7x41 multi_7x41_mod_52(clk,rst,matrix2_A[52],matrix2_B[52],mul_res2[52]);
multi_7x41 multi_7x41_mod_53(clk,rst,matrix2_A[53],matrix2_B[53],mul_res2[53]);
multi_7x41 multi_7x41_mod_54(clk,rst,matrix2_A[54],matrix2_B[54],mul_res2[54]);
multi_7x41 multi_7x41_mod_55(clk,rst,matrix2_A[55],matrix2_B[55],mul_res2[55]);
multi_7x41 multi_7x41_mod_56(clk,rst,matrix2_A[56],matrix2_B[56],mul_res2[56]);
multi_7x41 multi_7x41_mod_57(clk,rst,matrix2_A[57],matrix2_B[57],mul_res2[57]);
multi_7x41 multi_7x41_mod_58(clk,rst,matrix2_A[58],matrix2_B[58],mul_res2[58]);
multi_7x41 multi_7x41_mod_59(clk,rst,matrix2_A[59],matrix2_B[59],mul_res2[59]);
multi_7x41 multi_7x41_mod_60(clk,rst,matrix2_A[60],matrix2_B[60],mul_res2[60]);
multi_7x41 multi_7x41_mod_61(clk,rst,matrix2_A[61],matrix2_B[61],mul_res2[61]);
multi_7x41 multi_7x41_mod_62(clk,rst,matrix2_A[62],matrix2_B[62],mul_res2[62]);
multi_7x41 multi_7x41_mod_63(clk,rst,matrix2_A[63],matrix2_B[63],mul_res2[63]);
multi_7x41 multi_7x41_mod_64(clk,rst,matrix2_A[0],matrix2_B[64],mul_res2[64]);
multi_7x41 multi_7x41_mod_65(clk,rst,matrix2_A[1],matrix2_B[65],mul_res2[65]);
multi_7x41 multi_7x41_mod_66(clk,rst,matrix2_A[2],matrix2_B[66],mul_res2[66]);
multi_7x41 multi_7x41_mod_67(clk,rst,matrix2_A[3],matrix2_B[67],mul_res2[67]);
multi_7x41 multi_7x41_mod_68(clk,rst,matrix2_A[4],matrix2_B[68],mul_res2[68]);
multi_7x41 multi_7x41_mod_69(clk,rst,matrix2_A[5],matrix2_B[69],mul_res2[69]);
multi_7x41 multi_7x41_mod_70(clk,rst,matrix2_A[6],matrix2_B[70],mul_res2[70]);
multi_7x41 multi_7x41_mod_71(clk,rst,matrix2_A[7],matrix2_B[71],mul_res2[71]);
multi_7x41 multi_7x41_mod_72(clk,rst,matrix2_A[8],matrix2_B[72],mul_res2[72]);
multi_7x41 multi_7x41_mod_73(clk,rst,matrix2_A[9],matrix2_B[73],mul_res2[73]);
multi_7x41 multi_7x41_mod_74(clk,rst,matrix2_A[10],matrix2_B[74],mul_res2[74]);
multi_7x41 multi_7x41_mod_75(clk,rst,matrix2_A[11],matrix2_B[75],mul_res2[75]);
multi_7x41 multi_7x41_mod_76(clk,rst,matrix2_A[12],matrix2_B[76],mul_res2[76]);
multi_7x41 multi_7x41_mod_77(clk,rst,matrix2_A[13],matrix2_B[77],mul_res2[77]);
multi_7x41 multi_7x41_mod_78(clk,rst,matrix2_A[14],matrix2_B[78],mul_res2[78]);
multi_7x41 multi_7x41_mod_79(clk,rst,matrix2_A[15],matrix2_B[79],mul_res2[79]);
multi_7x41 multi_7x41_mod_80(clk,rst,matrix2_A[16],matrix2_B[80],mul_res2[80]);
multi_7x41 multi_7x41_mod_81(clk,rst,matrix2_A[17],matrix2_B[81],mul_res2[81]);
multi_7x41 multi_7x41_mod_82(clk,rst,matrix2_A[18],matrix2_B[82],mul_res2[82]);
multi_7x41 multi_7x41_mod_83(clk,rst,matrix2_A[19],matrix2_B[83],mul_res2[83]);
multi_7x41 multi_7x41_mod_84(clk,rst,matrix2_A[20],matrix2_B[84],mul_res2[84]);
multi_7x41 multi_7x41_mod_85(clk,rst,matrix2_A[21],matrix2_B[85],mul_res2[85]);
multi_7x41 multi_7x41_mod_86(clk,rst,matrix2_A[22],matrix2_B[86],mul_res2[86]);
multi_7x41 multi_7x41_mod_87(clk,rst,matrix2_A[23],matrix2_B[87],mul_res2[87]);
multi_7x41 multi_7x41_mod_88(clk,rst,matrix2_A[24],matrix2_B[88],mul_res2[88]);
multi_7x41 multi_7x41_mod_89(clk,rst,matrix2_A[25],matrix2_B[89],mul_res2[89]);
multi_7x41 multi_7x41_mod_90(clk,rst,matrix2_A[26],matrix2_B[90],mul_res2[90]);
multi_7x41 multi_7x41_mod_91(clk,rst,matrix2_A[27],matrix2_B[91],mul_res2[91]);
multi_7x41 multi_7x41_mod_92(clk,rst,matrix2_A[28],matrix2_B[92],mul_res2[92]);
multi_7x41 multi_7x41_mod_93(clk,rst,matrix2_A[29],matrix2_B[93],mul_res2[93]);
multi_7x41 multi_7x41_mod_94(clk,rst,matrix2_A[30],matrix2_B[94],mul_res2[94]);
multi_7x41 multi_7x41_mod_95(clk,rst,matrix2_A[31],matrix2_B[95],mul_res2[95]);
multi_7x41 multi_7x41_mod_96(clk,rst,matrix2_A[32],matrix2_B[96],mul_res2[96]);
multi_7x41 multi_7x41_mod_97(clk,rst,matrix2_A[33],matrix2_B[97],mul_res2[97]);
multi_7x41 multi_7x41_mod_98(clk,rst,matrix2_A[34],matrix2_B[98],mul_res2[98]);
multi_7x41 multi_7x41_mod_99(clk,rst,matrix2_A[35],matrix2_B[99],mul_res2[99]);
multi_7x41 multi_7x41_mod_100(clk,rst,matrix2_A[36],matrix2_B[100],mul_res2[100]);
multi_7x41 multi_7x41_mod_101(clk,rst,matrix2_A[37],matrix2_B[101],mul_res2[101]);
multi_7x41 multi_7x41_mod_102(clk,rst,matrix2_A[38],matrix2_B[102],mul_res2[102]);
multi_7x41 multi_7x41_mod_103(clk,rst,matrix2_A[39],matrix2_B[103],mul_res2[103]);
multi_7x41 multi_7x41_mod_104(clk,rst,matrix2_A[40],matrix2_B[104],mul_res2[104]);
multi_7x41 multi_7x41_mod_105(clk,rst,matrix2_A[41],matrix2_B[105],mul_res2[105]);
multi_7x41 multi_7x41_mod_106(clk,rst,matrix2_A[42],matrix2_B[106],mul_res2[106]);
multi_7x41 multi_7x41_mod_107(clk,rst,matrix2_A[43],matrix2_B[107],mul_res2[107]);
multi_7x41 multi_7x41_mod_108(clk,rst,matrix2_A[44],matrix2_B[108],mul_res2[108]);
multi_7x41 multi_7x41_mod_109(clk,rst,matrix2_A[45],matrix2_B[109],mul_res2[109]);
multi_7x41 multi_7x41_mod_110(clk,rst,matrix2_A[46],matrix2_B[110],mul_res2[110]);
multi_7x41 multi_7x41_mod_111(clk,rst,matrix2_A[47],matrix2_B[111],mul_res2[111]);
multi_7x41 multi_7x41_mod_112(clk,rst,matrix2_A[48],matrix2_B[112],mul_res2[112]);
multi_7x41 multi_7x41_mod_113(clk,rst,matrix2_A[49],matrix2_B[113],mul_res2[113]);
multi_7x41 multi_7x41_mod_114(clk,rst,matrix2_A[50],matrix2_B[114],mul_res2[114]);
multi_7x41 multi_7x41_mod_115(clk,rst,matrix2_A[51],matrix2_B[115],mul_res2[115]);
multi_7x41 multi_7x41_mod_116(clk,rst,matrix2_A[52],matrix2_B[116],mul_res2[116]);
multi_7x41 multi_7x41_mod_117(clk,rst,matrix2_A[53],matrix2_B[117],mul_res2[117]);
multi_7x41 multi_7x41_mod_118(clk,rst,matrix2_A[54],matrix2_B[118],mul_res2[118]);
multi_7x41 multi_7x41_mod_119(clk,rst,matrix2_A[55],matrix2_B[119],mul_res2[119]);
multi_7x41 multi_7x41_mod_120(clk,rst,matrix2_A[56],matrix2_B[120],mul_res2[120]);
multi_7x41 multi_7x41_mod_121(clk,rst,matrix2_A[57],matrix2_B[121],mul_res2[121]);
multi_7x41 multi_7x41_mod_122(clk,rst,matrix2_A[58],matrix2_B[122],mul_res2[122]);
multi_7x41 multi_7x41_mod_123(clk,rst,matrix2_A[59],matrix2_B[123],mul_res2[123]);
multi_7x41 multi_7x41_mod_124(clk,rst,matrix2_A[60],matrix2_B[124],mul_res2[124]);
multi_7x41 multi_7x41_mod_125(clk,rst,matrix2_A[61],matrix2_B[125],mul_res2[125]);
multi_7x41 multi_7x41_mod_126(clk,rst,matrix2_A[62],matrix2_B[126],mul_res2[126]);
multi_7x41 multi_7x41_mod_127(clk,rst,matrix2_A[63],matrix2_B[127],mul_res2[127]);
multi_7x41 multi_7x41_mod_128(clk,rst,matrix2_A[0],matrix2_B[128],mul_res2[128]);
multi_7x41 multi_7x41_mod_129(clk,rst,matrix2_A[1],matrix2_B[129],mul_res2[129]);
multi_7x41 multi_7x41_mod_130(clk,rst,matrix2_A[2],matrix2_B[130],mul_res2[130]);
multi_7x41 multi_7x41_mod_131(clk,rst,matrix2_A[3],matrix2_B[131],mul_res2[131]);
multi_7x41 multi_7x41_mod_132(clk,rst,matrix2_A[4],matrix2_B[132],mul_res2[132]);
multi_7x41 multi_7x41_mod_133(clk,rst,matrix2_A[5],matrix2_B[133],mul_res2[133]);
multi_7x41 multi_7x41_mod_134(clk,rst,matrix2_A[6],matrix2_B[134],mul_res2[134]);
multi_7x41 multi_7x41_mod_135(clk,rst,matrix2_A[7],matrix2_B[135],mul_res2[135]);
multi_7x41 multi_7x41_mod_136(clk,rst,matrix2_A[8],matrix2_B[136],mul_res2[136]);
multi_7x41 multi_7x41_mod_137(clk,rst,matrix2_A[9],matrix2_B[137],mul_res2[137]);
multi_7x41 multi_7x41_mod_138(clk,rst,matrix2_A[10],matrix2_B[138],mul_res2[138]);
multi_7x41 multi_7x41_mod_139(clk,rst,matrix2_A[11],matrix2_B[139],mul_res2[139]);
multi_7x41 multi_7x41_mod_140(clk,rst,matrix2_A[12],matrix2_B[140],mul_res2[140]);
multi_7x41 multi_7x41_mod_141(clk,rst,matrix2_A[13],matrix2_B[141],mul_res2[141]);
multi_7x41 multi_7x41_mod_142(clk,rst,matrix2_A[14],matrix2_B[142],mul_res2[142]);
multi_7x41 multi_7x41_mod_143(clk,rst,matrix2_A[15],matrix2_B[143],mul_res2[143]);
multi_7x41 multi_7x41_mod_144(clk,rst,matrix2_A[16],matrix2_B[144],mul_res2[144]);
multi_7x41 multi_7x41_mod_145(clk,rst,matrix2_A[17],matrix2_B[145],mul_res2[145]);
multi_7x41 multi_7x41_mod_146(clk,rst,matrix2_A[18],matrix2_B[146],mul_res2[146]);
multi_7x41 multi_7x41_mod_147(clk,rst,matrix2_A[19],matrix2_B[147],mul_res2[147]);
multi_7x41 multi_7x41_mod_148(clk,rst,matrix2_A[20],matrix2_B[148],mul_res2[148]);
multi_7x41 multi_7x41_mod_149(clk,rst,matrix2_A[21],matrix2_B[149],mul_res2[149]);
multi_7x41 multi_7x41_mod_150(clk,rst,matrix2_A[22],matrix2_B[150],mul_res2[150]);
multi_7x41 multi_7x41_mod_151(clk,rst,matrix2_A[23],matrix2_B[151],mul_res2[151]);
multi_7x41 multi_7x41_mod_152(clk,rst,matrix2_A[24],matrix2_B[152],mul_res2[152]);
multi_7x41 multi_7x41_mod_153(clk,rst,matrix2_A[25],matrix2_B[153],mul_res2[153]);
multi_7x41 multi_7x41_mod_154(clk,rst,matrix2_A[26],matrix2_B[154],mul_res2[154]);
multi_7x41 multi_7x41_mod_155(clk,rst,matrix2_A[27],matrix2_B[155],mul_res2[155]);
multi_7x41 multi_7x41_mod_156(clk,rst,matrix2_A[28],matrix2_B[156],mul_res2[156]);
multi_7x41 multi_7x41_mod_157(clk,rst,matrix2_A[29],matrix2_B[157],mul_res2[157]);
multi_7x41 multi_7x41_mod_158(clk,rst,matrix2_A[30],matrix2_B[158],mul_res2[158]);
multi_7x41 multi_7x41_mod_159(clk,rst,matrix2_A[31],matrix2_B[159],mul_res2[159]);
multi_7x41 multi_7x41_mod_160(clk,rst,matrix2_A[32],matrix2_B[160],mul_res2[160]);
multi_7x41 multi_7x41_mod_161(clk,rst,matrix2_A[33],matrix2_B[161],mul_res2[161]);
multi_7x41 multi_7x41_mod_162(clk,rst,matrix2_A[34],matrix2_B[162],mul_res2[162]);
multi_7x41 multi_7x41_mod_163(clk,rst,matrix2_A[35],matrix2_B[163],mul_res2[163]);
multi_7x41 multi_7x41_mod_164(clk,rst,matrix2_A[36],matrix2_B[164],mul_res2[164]);
multi_7x41 multi_7x41_mod_165(clk,rst,matrix2_A[37],matrix2_B[165],mul_res2[165]);
multi_7x41 multi_7x41_mod_166(clk,rst,matrix2_A[38],matrix2_B[166],mul_res2[166]);
multi_7x41 multi_7x41_mod_167(clk,rst,matrix2_A[39],matrix2_B[167],mul_res2[167]);
multi_7x41 multi_7x41_mod_168(clk,rst,matrix2_A[40],matrix2_B[168],mul_res2[168]);
multi_7x41 multi_7x41_mod_169(clk,rst,matrix2_A[41],matrix2_B[169],mul_res2[169]);
multi_7x41 multi_7x41_mod_170(clk,rst,matrix2_A[42],matrix2_B[170],mul_res2[170]);
multi_7x41 multi_7x41_mod_171(clk,rst,matrix2_A[43],matrix2_B[171],mul_res2[171]);
multi_7x41 multi_7x41_mod_172(clk,rst,matrix2_A[44],matrix2_B[172],mul_res2[172]);
multi_7x41 multi_7x41_mod_173(clk,rst,matrix2_A[45],matrix2_B[173],mul_res2[173]);
multi_7x41 multi_7x41_mod_174(clk,rst,matrix2_A[46],matrix2_B[174],mul_res2[174]);
multi_7x41 multi_7x41_mod_175(clk,rst,matrix2_A[47],matrix2_B[175],mul_res2[175]);
multi_7x41 multi_7x41_mod_176(clk,rst,matrix2_A[48],matrix2_B[176],mul_res2[176]);
multi_7x41 multi_7x41_mod_177(clk,rst,matrix2_A[49],matrix2_B[177],mul_res2[177]);
multi_7x41 multi_7x41_mod_178(clk,rst,matrix2_A[50],matrix2_B[178],mul_res2[178]);
multi_7x41 multi_7x41_mod_179(clk,rst,matrix2_A[51],matrix2_B[179],mul_res2[179]);
multi_7x41 multi_7x41_mod_180(clk,rst,matrix2_A[52],matrix2_B[180],mul_res2[180]);
multi_7x41 multi_7x41_mod_181(clk,rst,matrix2_A[53],matrix2_B[181],mul_res2[181]);
multi_7x41 multi_7x41_mod_182(clk,rst,matrix2_A[54],matrix2_B[182],mul_res2[182]);
multi_7x41 multi_7x41_mod_183(clk,rst,matrix2_A[55],matrix2_B[183],mul_res2[183]);
multi_7x41 multi_7x41_mod_184(clk,rst,matrix2_A[56],matrix2_B[184],mul_res2[184]);
multi_7x41 multi_7x41_mod_185(clk,rst,matrix2_A[57],matrix2_B[185],mul_res2[185]);
multi_7x41 multi_7x41_mod_186(clk,rst,matrix2_A[58],matrix2_B[186],mul_res2[186]);
multi_7x41 multi_7x41_mod_187(clk,rst,matrix2_A[59],matrix2_B[187],mul_res2[187]);
multi_7x41 multi_7x41_mod_188(clk,rst,matrix2_A[60],matrix2_B[188],mul_res2[188]);
multi_7x41 multi_7x41_mod_189(clk,rst,matrix2_A[61],matrix2_B[189],mul_res2[189]);
multi_7x41 multi_7x41_mod_190(clk,rst,matrix2_A[62],matrix2_B[190],mul_res2[190]);
multi_7x41 multi_7x41_mod_191(clk,rst,matrix2_A[63],matrix2_B[191],mul_res2[191]);
multi_7x41 multi_7x41_mod_192(clk,rst,matrix2_A[0],matrix2_B[192],mul_res2[192]);
multi_7x41 multi_7x41_mod_193(clk,rst,matrix2_A[1],matrix2_B[193],mul_res2[193]);
multi_7x41 multi_7x41_mod_194(clk,rst,matrix2_A[2],matrix2_B[194],mul_res2[194]);
multi_7x41 multi_7x41_mod_195(clk,rst,matrix2_A[3],matrix2_B[195],mul_res2[195]);
multi_7x41 multi_7x41_mod_196(clk,rst,matrix2_A[4],matrix2_B[196],mul_res2[196]);
multi_7x41 multi_7x41_mod_197(clk,rst,matrix2_A[5],matrix2_B[197],mul_res2[197]);
multi_7x41 multi_7x41_mod_198(clk,rst,matrix2_A[6],matrix2_B[198],mul_res2[198]);
multi_7x41 multi_7x41_mod_199(clk,rst,matrix2_A[7],matrix2_B[199],mul_res2[199]);
multi_7x41 multi_7x41_mod_200(clk,rst,matrix2_A[8],matrix2_B[200],mul_res2[200]);
multi_7x41 multi_7x41_mod_201(clk,rst,matrix2_A[9],matrix2_B[201],mul_res2[201]);
multi_7x41 multi_7x41_mod_202(clk,rst,matrix2_A[10],matrix2_B[202],mul_res2[202]);
multi_7x41 multi_7x41_mod_203(clk,rst,matrix2_A[11],matrix2_B[203],mul_res2[203]);
multi_7x41 multi_7x41_mod_204(clk,rst,matrix2_A[12],matrix2_B[204],mul_res2[204]);
multi_7x41 multi_7x41_mod_205(clk,rst,matrix2_A[13],matrix2_B[205],mul_res2[205]);
multi_7x41 multi_7x41_mod_206(clk,rst,matrix2_A[14],matrix2_B[206],mul_res2[206]);
multi_7x41 multi_7x41_mod_207(clk,rst,matrix2_A[15],matrix2_B[207],mul_res2[207]);
multi_7x41 multi_7x41_mod_208(clk,rst,matrix2_A[16],matrix2_B[208],mul_res2[208]);
multi_7x41 multi_7x41_mod_209(clk,rst,matrix2_A[17],matrix2_B[209],mul_res2[209]);
multi_7x41 multi_7x41_mod_210(clk,rst,matrix2_A[18],matrix2_B[210],mul_res2[210]);
multi_7x41 multi_7x41_mod_211(clk,rst,matrix2_A[19],matrix2_B[211],mul_res2[211]);
multi_7x41 multi_7x41_mod_212(clk,rst,matrix2_A[20],matrix2_B[212],mul_res2[212]);
multi_7x41 multi_7x41_mod_213(clk,rst,matrix2_A[21],matrix2_B[213],mul_res2[213]);
multi_7x41 multi_7x41_mod_214(clk,rst,matrix2_A[22],matrix2_B[214],mul_res2[214]);
multi_7x41 multi_7x41_mod_215(clk,rst,matrix2_A[23],matrix2_B[215],mul_res2[215]);
multi_7x41 multi_7x41_mod_216(clk,rst,matrix2_A[24],matrix2_B[216],mul_res2[216]);
multi_7x41 multi_7x41_mod_217(clk,rst,matrix2_A[25],matrix2_B[217],mul_res2[217]);
multi_7x41 multi_7x41_mod_218(clk,rst,matrix2_A[26],matrix2_B[218],mul_res2[218]);
multi_7x41 multi_7x41_mod_219(clk,rst,matrix2_A[27],matrix2_B[219],mul_res2[219]);
multi_7x41 multi_7x41_mod_220(clk,rst,matrix2_A[28],matrix2_B[220],mul_res2[220]);
multi_7x41 multi_7x41_mod_221(clk,rst,matrix2_A[29],matrix2_B[221],mul_res2[221]);
multi_7x41 multi_7x41_mod_222(clk,rst,matrix2_A[30],matrix2_B[222],mul_res2[222]);
multi_7x41 multi_7x41_mod_223(clk,rst,matrix2_A[31],matrix2_B[223],mul_res2[223]);
multi_7x41 multi_7x41_mod_224(clk,rst,matrix2_A[32],matrix2_B[224],mul_res2[224]);
multi_7x41 multi_7x41_mod_225(clk,rst,matrix2_A[33],matrix2_B[225],mul_res2[225]);
multi_7x41 multi_7x41_mod_226(clk,rst,matrix2_A[34],matrix2_B[226],mul_res2[226]);
multi_7x41 multi_7x41_mod_227(clk,rst,matrix2_A[35],matrix2_B[227],mul_res2[227]);
multi_7x41 multi_7x41_mod_228(clk,rst,matrix2_A[36],matrix2_B[228],mul_res2[228]);
multi_7x41 multi_7x41_mod_229(clk,rst,matrix2_A[37],matrix2_B[229],mul_res2[229]);
multi_7x41 multi_7x41_mod_230(clk,rst,matrix2_A[38],matrix2_B[230],mul_res2[230]);
multi_7x41 multi_7x41_mod_231(clk,rst,matrix2_A[39],matrix2_B[231],mul_res2[231]);
multi_7x41 multi_7x41_mod_232(clk,rst,matrix2_A[40],matrix2_B[232],mul_res2[232]);
multi_7x41 multi_7x41_mod_233(clk,rst,matrix2_A[41],matrix2_B[233],mul_res2[233]);
multi_7x41 multi_7x41_mod_234(clk,rst,matrix2_A[42],matrix2_B[234],mul_res2[234]);
multi_7x41 multi_7x41_mod_235(clk,rst,matrix2_A[43],matrix2_B[235],mul_res2[235]);
multi_7x41 multi_7x41_mod_236(clk,rst,matrix2_A[44],matrix2_B[236],mul_res2[236]);
multi_7x41 multi_7x41_mod_237(clk,rst,matrix2_A[45],matrix2_B[237],mul_res2[237]);
multi_7x41 multi_7x41_mod_238(clk,rst,matrix2_A[46],matrix2_B[238],mul_res2[238]);
multi_7x41 multi_7x41_mod_239(clk,rst,matrix2_A[47],matrix2_B[239],mul_res2[239]);
multi_7x41 multi_7x41_mod_240(clk,rst,matrix2_A[48],matrix2_B[240],mul_res2[240]);
multi_7x41 multi_7x41_mod_241(clk,rst,matrix2_A[49],matrix2_B[241],mul_res2[241]);
multi_7x41 multi_7x41_mod_242(clk,rst,matrix2_A[50],matrix2_B[242],mul_res2[242]);
multi_7x41 multi_7x41_mod_243(clk,rst,matrix2_A[51],matrix2_B[243],mul_res2[243]);
multi_7x41 multi_7x41_mod_244(clk,rst,matrix2_A[52],matrix2_B[244],mul_res2[244]);
multi_7x41 multi_7x41_mod_245(clk,rst,matrix2_A[53],matrix2_B[245],mul_res2[245]);
multi_7x41 multi_7x41_mod_246(clk,rst,matrix2_A[54],matrix2_B[246],mul_res2[246]);
multi_7x41 multi_7x41_mod_247(clk,rst,matrix2_A[55],matrix2_B[247],mul_res2[247]);
multi_7x41 multi_7x41_mod_248(clk,rst,matrix2_A[56],matrix2_B[248],mul_res2[248]);
multi_7x41 multi_7x41_mod_249(clk,rst,matrix2_A[57],matrix2_B[249],mul_res2[249]);
multi_7x41 multi_7x41_mod_250(clk,rst,matrix2_A[58],matrix2_B[250],mul_res2[250]);
multi_7x41 multi_7x41_mod_251(clk,rst,matrix2_A[59],matrix2_B[251],mul_res2[251]);
multi_7x41 multi_7x41_mod_252(clk,rst,matrix2_A[60],matrix2_B[252],mul_res2[252]);
multi_7x41 multi_7x41_mod_253(clk,rst,matrix2_A[61],matrix2_B[253],mul_res2[253]);
multi_7x41 multi_7x41_mod_254(clk,rst,matrix2_A[62],matrix2_B[254],mul_res2[254]);
multi_7x41 multi_7x41_mod_255(clk,rst,matrix2_A[63],matrix2_B[255],mul_res2[255]);
multi_7x41 multi_7x41_mod_256(clk,rst,matrix2_A[0],matrix2_B[256],mul_res2[256]);
multi_7x41 multi_7x41_mod_257(clk,rst,matrix2_A[1],matrix2_B[257],mul_res2[257]);
multi_7x41 multi_7x41_mod_258(clk,rst,matrix2_A[2],matrix2_B[258],mul_res2[258]);
multi_7x41 multi_7x41_mod_259(clk,rst,matrix2_A[3],matrix2_B[259],mul_res2[259]);
multi_7x41 multi_7x41_mod_260(clk,rst,matrix2_A[4],matrix2_B[260],mul_res2[260]);
multi_7x41 multi_7x41_mod_261(clk,rst,matrix2_A[5],matrix2_B[261],mul_res2[261]);
multi_7x41 multi_7x41_mod_262(clk,rst,matrix2_A[6],matrix2_B[262],mul_res2[262]);
multi_7x41 multi_7x41_mod_263(clk,rst,matrix2_A[7],matrix2_B[263],mul_res2[263]);
multi_7x41 multi_7x41_mod_264(clk,rst,matrix2_A[8],matrix2_B[264],mul_res2[264]);
multi_7x41 multi_7x41_mod_265(clk,rst,matrix2_A[9],matrix2_B[265],mul_res2[265]);
multi_7x41 multi_7x41_mod_266(clk,rst,matrix2_A[10],matrix2_B[266],mul_res2[266]);
multi_7x41 multi_7x41_mod_267(clk,rst,matrix2_A[11],matrix2_B[267],mul_res2[267]);
multi_7x41 multi_7x41_mod_268(clk,rst,matrix2_A[12],matrix2_B[268],mul_res2[268]);
multi_7x41 multi_7x41_mod_269(clk,rst,matrix2_A[13],matrix2_B[269],mul_res2[269]);
multi_7x41 multi_7x41_mod_270(clk,rst,matrix2_A[14],matrix2_B[270],mul_res2[270]);
multi_7x41 multi_7x41_mod_271(clk,rst,matrix2_A[15],matrix2_B[271],mul_res2[271]);
multi_7x41 multi_7x41_mod_272(clk,rst,matrix2_A[16],matrix2_B[272],mul_res2[272]);
multi_7x41 multi_7x41_mod_273(clk,rst,matrix2_A[17],matrix2_B[273],mul_res2[273]);
multi_7x41 multi_7x41_mod_274(clk,rst,matrix2_A[18],matrix2_B[274],mul_res2[274]);
multi_7x41 multi_7x41_mod_275(clk,rst,matrix2_A[19],matrix2_B[275],mul_res2[275]);
multi_7x41 multi_7x41_mod_276(clk,rst,matrix2_A[20],matrix2_B[276],mul_res2[276]);
multi_7x41 multi_7x41_mod_277(clk,rst,matrix2_A[21],matrix2_B[277],mul_res2[277]);
multi_7x41 multi_7x41_mod_278(clk,rst,matrix2_A[22],matrix2_B[278],mul_res2[278]);
multi_7x41 multi_7x41_mod_279(clk,rst,matrix2_A[23],matrix2_B[279],mul_res2[279]);
multi_7x41 multi_7x41_mod_280(clk,rst,matrix2_A[24],matrix2_B[280],mul_res2[280]);
multi_7x41 multi_7x41_mod_281(clk,rst,matrix2_A[25],matrix2_B[281],mul_res2[281]);
multi_7x41 multi_7x41_mod_282(clk,rst,matrix2_A[26],matrix2_B[282],mul_res2[282]);
multi_7x41 multi_7x41_mod_283(clk,rst,matrix2_A[27],matrix2_B[283],mul_res2[283]);
multi_7x41 multi_7x41_mod_284(clk,rst,matrix2_A[28],matrix2_B[284],mul_res2[284]);
multi_7x41 multi_7x41_mod_285(clk,rst,matrix2_A[29],matrix2_B[285],mul_res2[285]);
multi_7x41 multi_7x41_mod_286(clk,rst,matrix2_A[30],matrix2_B[286],mul_res2[286]);
multi_7x41 multi_7x41_mod_287(clk,rst,matrix2_A[31],matrix2_B[287],mul_res2[287]);
multi_7x41 multi_7x41_mod_288(clk,rst,matrix2_A[32],matrix2_B[288],mul_res2[288]);
multi_7x41 multi_7x41_mod_289(clk,rst,matrix2_A[33],matrix2_B[289],mul_res2[289]);
multi_7x41 multi_7x41_mod_290(clk,rst,matrix2_A[34],matrix2_B[290],mul_res2[290]);
multi_7x41 multi_7x41_mod_291(clk,rst,matrix2_A[35],matrix2_B[291],mul_res2[291]);
multi_7x41 multi_7x41_mod_292(clk,rst,matrix2_A[36],matrix2_B[292],mul_res2[292]);
multi_7x41 multi_7x41_mod_293(clk,rst,matrix2_A[37],matrix2_B[293],mul_res2[293]);
multi_7x41 multi_7x41_mod_294(clk,rst,matrix2_A[38],matrix2_B[294],mul_res2[294]);
multi_7x41 multi_7x41_mod_295(clk,rst,matrix2_A[39],matrix2_B[295],mul_res2[295]);
multi_7x41 multi_7x41_mod_296(clk,rst,matrix2_A[40],matrix2_B[296],mul_res2[296]);
multi_7x41 multi_7x41_mod_297(clk,rst,matrix2_A[41],matrix2_B[297],mul_res2[297]);
multi_7x41 multi_7x41_mod_298(clk,rst,matrix2_A[42],matrix2_B[298],mul_res2[298]);
multi_7x41 multi_7x41_mod_299(clk,rst,matrix2_A[43],matrix2_B[299],mul_res2[299]);
multi_7x41 multi_7x41_mod_300(clk,rst,matrix2_A[44],matrix2_B[300],mul_res2[300]);
multi_7x41 multi_7x41_mod_301(clk,rst,matrix2_A[45],matrix2_B[301],mul_res2[301]);
multi_7x41 multi_7x41_mod_302(clk,rst,matrix2_A[46],matrix2_B[302],mul_res2[302]);
multi_7x41 multi_7x41_mod_303(clk,rst,matrix2_A[47],matrix2_B[303],mul_res2[303]);
multi_7x41 multi_7x41_mod_304(clk,rst,matrix2_A[48],matrix2_B[304],mul_res2[304]);
multi_7x41 multi_7x41_mod_305(clk,rst,matrix2_A[49],matrix2_B[305],mul_res2[305]);
multi_7x41 multi_7x41_mod_306(clk,rst,matrix2_A[50],matrix2_B[306],mul_res2[306]);
multi_7x41 multi_7x41_mod_307(clk,rst,matrix2_A[51],matrix2_B[307],mul_res2[307]);
multi_7x41 multi_7x41_mod_308(clk,rst,matrix2_A[52],matrix2_B[308],mul_res2[308]);
multi_7x41 multi_7x41_mod_309(clk,rst,matrix2_A[53],matrix2_B[309],mul_res2[309]);
multi_7x41 multi_7x41_mod_310(clk,rst,matrix2_A[54],matrix2_B[310],mul_res2[310]);
multi_7x41 multi_7x41_mod_311(clk,rst,matrix2_A[55],matrix2_B[311],mul_res2[311]);
multi_7x41 multi_7x41_mod_312(clk,rst,matrix2_A[56],matrix2_B[312],mul_res2[312]);
multi_7x41 multi_7x41_mod_313(clk,rst,matrix2_A[57],matrix2_B[313],mul_res2[313]);
multi_7x41 multi_7x41_mod_314(clk,rst,matrix2_A[58],matrix2_B[314],mul_res2[314]);
multi_7x41 multi_7x41_mod_315(clk,rst,matrix2_A[59],matrix2_B[315],mul_res2[315]);
multi_7x41 multi_7x41_mod_316(clk,rst,matrix2_A[60],matrix2_B[316],mul_res2[316]);
multi_7x41 multi_7x41_mod_317(clk,rst,matrix2_A[61],matrix2_B[317],mul_res2[317]);
multi_7x41 multi_7x41_mod_318(clk,rst,matrix2_A[62],matrix2_B[318],mul_res2[318]);
multi_7x41 multi_7x41_mod_319(clk,rst,matrix2_A[63],matrix2_B[319],mul_res2[319]);
multi_7x41 multi_7x41_mod_320(clk,rst,matrix2_A[0],matrix2_B[320],mul_res2[320]);
multi_7x41 multi_7x41_mod_321(clk,rst,matrix2_A[1],matrix2_B[321],mul_res2[321]);
multi_7x41 multi_7x41_mod_322(clk,rst,matrix2_A[2],matrix2_B[322],mul_res2[322]);
multi_7x41 multi_7x41_mod_323(clk,rst,matrix2_A[3],matrix2_B[323],mul_res2[323]);
multi_7x41 multi_7x41_mod_324(clk,rst,matrix2_A[4],matrix2_B[324],mul_res2[324]);
multi_7x41 multi_7x41_mod_325(clk,rst,matrix2_A[5],matrix2_B[325],mul_res2[325]);
multi_7x41 multi_7x41_mod_326(clk,rst,matrix2_A[6],matrix2_B[326],mul_res2[326]);
multi_7x41 multi_7x41_mod_327(clk,rst,matrix2_A[7],matrix2_B[327],mul_res2[327]);
multi_7x41 multi_7x41_mod_328(clk,rst,matrix2_A[8],matrix2_B[328],mul_res2[328]);
multi_7x41 multi_7x41_mod_329(clk,rst,matrix2_A[9],matrix2_B[329],mul_res2[329]);
multi_7x41 multi_7x41_mod_330(clk,rst,matrix2_A[10],matrix2_B[330],mul_res2[330]);
multi_7x41 multi_7x41_mod_331(clk,rst,matrix2_A[11],matrix2_B[331],mul_res2[331]);
multi_7x41 multi_7x41_mod_332(clk,rst,matrix2_A[12],matrix2_B[332],mul_res2[332]);
multi_7x41 multi_7x41_mod_333(clk,rst,matrix2_A[13],matrix2_B[333],mul_res2[333]);
multi_7x41 multi_7x41_mod_334(clk,rst,matrix2_A[14],matrix2_B[334],mul_res2[334]);
multi_7x41 multi_7x41_mod_335(clk,rst,matrix2_A[15],matrix2_B[335],mul_res2[335]);
multi_7x41 multi_7x41_mod_336(clk,rst,matrix2_A[16],matrix2_B[336],mul_res2[336]);
multi_7x41 multi_7x41_mod_337(clk,rst,matrix2_A[17],matrix2_B[337],mul_res2[337]);
multi_7x41 multi_7x41_mod_338(clk,rst,matrix2_A[18],matrix2_B[338],mul_res2[338]);
multi_7x41 multi_7x41_mod_339(clk,rst,matrix2_A[19],matrix2_B[339],mul_res2[339]);
multi_7x41 multi_7x41_mod_340(clk,rst,matrix2_A[20],matrix2_B[340],mul_res2[340]);
multi_7x41 multi_7x41_mod_341(clk,rst,matrix2_A[21],matrix2_B[341],mul_res2[341]);
multi_7x41 multi_7x41_mod_342(clk,rst,matrix2_A[22],matrix2_B[342],mul_res2[342]);
multi_7x41 multi_7x41_mod_343(clk,rst,matrix2_A[23],matrix2_B[343],mul_res2[343]);
multi_7x41 multi_7x41_mod_344(clk,rst,matrix2_A[24],matrix2_B[344],mul_res2[344]);
multi_7x41 multi_7x41_mod_345(clk,rst,matrix2_A[25],matrix2_B[345],mul_res2[345]);
multi_7x41 multi_7x41_mod_346(clk,rst,matrix2_A[26],matrix2_B[346],mul_res2[346]);
multi_7x41 multi_7x41_mod_347(clk,rst,matrix2_A[27],matrix2_B[347],mul_res2[347]);
multi_7x41 multi_7x41_mod_348(clk,rst,matrix2_A[28],matrix2_B[348],mul_res2[348]);
multi_7x41 multi_7x41_mod_349(clk,rst,matrix2_A[29],matrix2_B[349],mul_res2[349]);
multi_7x41 multi_7x41_mod_350(clk,rst,matrix2_A[30],matrix2_B[350],mul_res2[350]);
multi_7x41 multi_7x41_mod_351(clk,rst,matrix2_A[31],matrix2_B[351],mul_res2[351]);
multi_7x41 multi_7x41_mod_352(clk,rst,matrix2_A[32],matrix2_B[352],mul_res2[352]);
multi_7x41 multi_7x41_mod_353(clk,rst,matrix2_A[33],matrix2_B[353],mul_res2[353]);
multi_7x41 multi_7x41_mod_354(clk,rst,matrix2_A[34],matrix2_B[354],mul_res2[354]);
multi_7x41 multi_7x41_mod_355(clk,rst,matrix2_A[35],matrix2_B[355],mul_res2[355]);
multi_7x41 multi_7x41_mod_356(clk,rst,matrix2_A[36],matrix2_B[356],mul_res2[356]);
multi_7x41 multi_7x41_mod_357(clk,rst,matrix2_A[37],matrix2_B[357],mul_res2[357]);
multi_7x41 multi_7x41_mod_358(clk,rst,matrix2_A[38],matrix2_B[358],mul_res2[358]);
multi_7x41 multi_7x41_mod_359(clk,rst,matrix2_A[39],matrix2_B[359],mul_res2[359]);
multi_7x41 multi_7x41_mod_360(clk,rst,matrix2_A[40],matrix2_B[360],mul_res2[360]);
multi_7x41 multi_7x41_mod_361(clk,rst,matrix2_A[41],matrix2_B[361],mul_res2[361]);
multi_7x41 multi_7x41_mod_362(clk,rst,matrix2_A[42],matrix2_B[362],mul_res2[362]);
multi_7x41 multi_7x41_mod_363(clk,rst,matrix2_A[43],matrix2_B[363],mul_res2[363]);
multi_7x41 multi_7x41_mod_364(clk,rst,matrix2_A[44],matrix2_B[364],mul_res2[364]);
multi_7x41 multi_7x41_mod_365(clk,rst,matrix2_A[45],matrix2_B[365],mul_res2[365]);
multi_7x41 multi_7x41_mod_366(clk,rst,matrix2_A[46],matrix2_B[366],mul_res2[366]);
multi_7x41 multi_7x41_mod_367(clk,rst,matrix2_A[47],matrix2_B[367],mul_res2[367]);
multi_7x41 multi_7x41_mod_368(clk,rst,matrix2_A[48],matrix2_B[368],mul_res2[368]);
multi_7x41 multi_7x41_mod_369(clk,rst,matrix2_A[49],matrix2_B[369],mul_res2[369]);
multi_7x41 multi_7x41_mod_370(clk,rst,matrix2_A[50],matrix2_B[370],mul_res2[370]);
multi_7x41 multi_7x41_mod_371(clk,rst,matrix2_A[51],matrix2_B[371],mul_res2[371]);
multi_7x41 multi_7x41_mod_372(clk,rst,matrix2_A[52],matrix2_B[372],mul_res2[372]);
multi_7x41 multi_7x41_mod_373(clk,rst,matrix2_A[53],matrix2_B[373],mul_res2[373]);
multi_7x41 multi_7x41_mod_374(clk,rst,matrix2_A[54],matrix2_B[374],mul_res2[374]);
multi_7x41 multi_7x41_mod_375(clk,rst,matrix2_A[55],matrix2_B[375],mul_res2[375]);
multi_7x41 multi_7x41_mod_376(clk,rst,matrix2_A[56],matrix2_B[376],mul_res2[376]);
multi_7x41 multi_7x41_mod_377(clk,rst,matrix2_A[57],matrix2_B[377],mul_res2[377]);
multi_7x41 multi_7x41_mod_378(clk,rst,matrix2_A[58],matrix2_B[378],mul_res2[378]);
multi_7x41 multi_7x41_mod_379(clk,rst,matrix2_A[59],matrix2_B[379],mul_res2[379]);
multi_7x41 multi_7x41_mod_380(clk,rst,matrix2_A[60],matrix2_B[380],mul_res2[380]);
multi_7x41 multi_7x41_mod_381(clk,rst,matrix2_A[61],matrix2_B[381],mul_res2[381]);
multi_7x41 multi_7x41_mod_382(clk,rst,matrix2_A[62],matrix2_B[382],mul_res2[382]);
multi_7x41 multi_7x41_mod_383(clk,rst,matrix2_A[63],matrix2_B[383],mul_res2[383]);
multi_7x41 multi_7x41_mod_384(clk,rst,matrix2_A[0],matrix2_B[384],mul_res2[384]);
multi_7x41 multi_7x41_mod_385(clk,rst,matrix2_A[1],matrix2_B[385],mul_res2[385]);
multi_7x41 multi_7x41_mod_386(clk,rst,matrix2_A[2],matrix2_B[386],mul_res2[386]);
multi_7x41 multi_7x41_mod_387(clk,rst,matrix2_A[3],matrix2_B[387],mul_res2[387]);
multi_7x41 multi_7x41_mod_388(clk,rst,matrix2_A[4],matrix2_B[388],mul_res2[388]);
multi_7x41 multi_7x41_mod_389(clk,rst,matrix2_A[5],matrix2_B[389],mul_res2[389]);
multi_7x41 multi_7x41_mod_390(clk,rst,matrix2_A[6],matrix2_B[390],mul_res2[390]);
multi_7x41 multi_7x41_mod_391(clk,rst,matrix2_A[7],matrix2_B[391],mul_res2[391]);
multi_7x41 multi_7x41_mod_392(clk,rst,matrix2_A[8],matrix2_B[392],mul_res2[392]);
multi_7x41 multi_7x41_mod_393(clk,rst,matrix2_A[9],matrix2_B[393],mul_res2[393]);
multi_7x41 multi_7x41_mod_394(clk,rst,matrix2_A[10],matrix2_B[394],mul_res2[394]);
multi_7x41 multi_7x41_mod_395(clk,rst,matrix2_A[11],matrix2_B[395],mul_res2[395]);
multi_7x41 multi_7x41_mod_396(clk,rst,matrix2_A[12],matrix2_B[396],mul_res2[396]);
multi_7x41 multi_7x41_mod_397(clk,rst,matrix2_A[13],matrix2_B[397],mul_res2[397]);
multi_7x41 multi_7x41_mod_398(clk,rst,matrix2_A[14],matrix2_B[398],mul_res2[398]);
multi_7x41 multi_7x41_mod_399(clk,rst,matrix2_A[15],matrix2_B[399],mul_res2[399]);
multi_7x41 multi_7x41_mod_400(clk,rst,matrix2_A[16],matrix2_B[400],mul_res2[400]);
multi_7x41 multi_7x41_mod_401(clk,rst,matrix2_A[17],matrix2_B[401],mul_res2[401]);
multi_7x41 multi_7x41_mod_402(clk,rst,matrix2_A[18],matrix2_B[402],mul_res2[402]);
multi_7x41 multi_7x41_mod_403(clk,rst,matrix2_A[19],matrix2_B[403],mul_res2[403]);
multi_7x41 multi_7x41_mod_404(clk,rst,matrix2_A[20],matrix2_B[404],mul_res2[404]);
multi_7x41 multi_7x41_mod_405(clk,rst,matrix2_A[21],matrix2_B[405],mul_res2[405]);
multi_7x41 multi_7x41_mod_406(clk,rst,matrix2_A[22],matrix2_B[406],mul_res2[406]);
multi_7x41 multi_7x41_mod_407(clk,rst,matrix2_A[23],matrix2_B[407],mul_res2[407]);
multi_7x41 multi_7x41_mod_408(clk,rst,matrix2_A[24],matrix2_B[408],mul_res2[408]);
multi_7x41 multi_7x41_mod_409(clk,rst,matrix2_A[25],matrix2_B[409],mul_res2[409]);
multi_7x41 multi_7x41_mod_410(clk,rst,matrix2_A[26],matrix2_B[410],mul_res2[410]);
multi_7x41 multi_7x41_mod_411(clk,rst,matrix2_A[27],matrix2_B[411],mul_res2[411]);
multi_7x41 multi_7x41_mod_412(clk,rst,matrix2_A[28],matrix2_B[412],mul_res2[412]);
multi_7x41 multi_7x41_mod_413(clk,rst,matrix2_A[29],matrix2_B[413],mul_res2[413]);
multi_7x41 multi_7x41_mod_414(clk,rst,matrix2_A[30],matrix2_B[414],mul_res2[414]);
multi_7x41 multi_7x41_mod_415(clk,rst,matrix2_A[31],matrix2_B[415],mul_res2[415]);
multi_7x41 multi_7x41_mod_416(clk,rst,matrix2_A[32],matrix2_B[416],mul_res2[416]);
multi_7x41 multi_7x41_mod_417(clk,rst,matrix2_A[33],matrix2_B[417],mul_res2[417]);
multi_7x41 multi_7x41_mod_418(clk,rst,matrix2_A[34],matrix2_B[418],mul_res2[418]);
multi_7x41 multi_7x41_mod_419(clk,rst,matrix2_A[35],matrix2_B[419],mul_res2[419]);
multi_7x41 multi_7x41_mod_420(clk,rst,matrix2_A[36],matrix2_B[420],mul_res2[420]);
multi_7x41 multi_7x41_mod_421(clk,rst,matrix2_A[37],matrix2_B[421],mul_res2[421]);
multi_7x41 multi_7x41_mod_422(clk,rst,matrix2_A[38],matrix2_B[422],mul_res2[422]);
multi_7x41 multi_7x41_mod_423(clk,rst,matrix2_A[39],matrix2_B[423],mul_res2[423]);
multi_7x41 multi_7x41_mod_424(clk,rst,matrix2_A[40],matrix2_B[424],mul_res2[424]);
multi_7x41 multi_7x41_mod_425(clk,rst,matrix2_A[41],matrix2_B[425],mul_res2[425]);
multi_7x41 multi_7x41_mod_426(clk,rst,matrix2_A[42],matrix2_B[426],mul_res2[426]);
multi_7x41 multi_7x41_mod_427(clk,rst,matrix2_A[43],matrix2_B[427],mul_res2[427]);
multi_7x41 multi_7x41_mod_428(clk,rst,matrix2_A[44],matrix2_B[428],mul_res2[428]);
multi_7x41 multi_7x41_mod_429(clk,rst,matrix2_A[45],matrix2_B[429],mul_res2[429]);
multi_7x41 multi_7x41_mod_430(clk,rst,matrix2_A[46],matrix2_B[430],mul_res2[430]);
multi_7x41 multi_7x41_mod_431(clk,rst,matrix2_A[47],matrix2_B[431],mul_res2[431]);
multi_7x41 multi_7x41_mod_432(clk,rst,matrix2_A[48],matrix2_B[432],mul_res2[432]);
multi_7x41 multi_7x41_mod_433(clk,rst,matrix2_A[49],matrix2_B[433],mul_res2[433]);
multi_7x41 multi_7x41_mod_434(clk,rst,matrix2_A[50],matrix2_B[434],mul_res2[434]);
multi_7x41 multi_7x41_mod_435(clk,rst,matrix2_A[51],matrix2_B[435],mul_res2[435]);
multi_7x41 multi_7x41_mod_436(clk,rst,matrix2_A[52],matrix2_B[436],mul_res2[436]);
multi_7x41 multi_7x41_mod_437(clk,rst,matrix2_A[53],matrix2_B[437],mul_res2[437]);
multi_7x41 multi_7x41_mod_438(clk,rst,matrix2_A[54],matrix2_B[438],mul_res2[438]);
multi_7x41 multi_7x41_mod_439(clk,rst,matrix2_A[55],matrix2_B[439],mul_res2[439]);
multi_7x41 multi_7x41_mod_440(clk,rst,matrix2_A[56],matrix2_B[440],mul_res2[440]);
multi_7x41 multi_7x41_mod_441(clk,rst,matrix2_A[57],matrix2_B[441],mul_res2[441]);
multi_7x41 multi_7x41_mod_442(clk,rst,matrix2_A[58],matrix2_B[442],mul_res2[442]);
multi_7x41 multi_7x41_mod_443(clk,rst,matrix2_A[59],matrix2_B[443],mul_res2[443]);
multi_7x41 multi_7x41_mod_444(clk,rst,matrix2_A[60],matrix2_B[444],mul_res2[444]);
multi_7x41 multi_7x41_mod_445(clk,rst,matrix2_A[61],matrix2_B[445],mul_res2[445]);
multi_7x41 multi_7x41_mod_446(clk,rst,matrix2_A[62],matrix2_B[446],mul_res2[446]);
multi_7x41 multi_7x41_mod_447(clk,rst,matrix2_A[63],matrix2_B[447],mul_res2[447]);
multi_7x41 multi_7x41_mod_448(clk,rst,matrix2_A[0],matrix2_B[448],mul_res2[448]);
multi_7x41 multi_7x41_mod_449(clk,rst,matrix2_A[1],matrix2_B[449],mul_res2[449]);
multi_7x41 multi_7x41_mod_450(clk,rst,matrix2_A[2],matrix2_B[450],mul_res2[450]);
multi_7x41 multi_7x41_mod_451(clk,rst,matrix2_A[3],matrix2_B[451],mul_res2[451]);
multi_7x41 multi_7x41_mod_452(clk,rst,matrix2_A[4],matrix2_B[452],mul_res2[452]);
multi_7x41 multi_7x41_mod_453(clk,rst,matrix2_A[5],matrix2_B[453],mul_res2[453]);
multi_7x41 multi_7x41_mod_454(clk,rst,matrix2_A[6],matrix2_B[454],mul_res2[454]);
multi_7x41 multi_7x41_mod_455(clk,rst,matrix2_A[7],matrix2_B[455],mul_res2[455]);
multi_7x41 multi_7x41_mod_456(clk,rst,matrix2_A[8],matrix2_B[456],mul_res2[456]);
multi_7x41 multi_7x41_mod_457(clk,rst,matrix2_A[9],matrix2_B[457],mul_res2[457]);
multi_7x41 multi_7x41_mod_458(clk,rst,matrix2_A[10],matrix2_B[458],mul_res2[458]);
multi_7x41 multi_7x41_mod_459(clk,rst,matrix2_A[11],matrix2_B[459],mul_res2[459]);
multi_7x41 multi_7x41_mod_460(clk,rst,matrix2_A[12],matrix2_B[460],mul_res2[460]);
multi_7x41 multi_7x41_mod_461(clk,rst,matrix2_A[13],matrix2_B[461],mul_res2[461]);
multi_7x41 multi_7x41_mod_462(clk,rst,matrix2_A[14],matrix2_B[462],mul_res2[462]);
multi_7x41 multi_7x41_mod_463(clk,rst,matrix2_A[15],matrix2_B[463],mul_res2[463]);
multi_7x41 multi_7x41_mod_464(clk,rst,matrix2_A[16],matrix2_B[464],mul_res2[464]);
multi_7x41 multi_7x41_mod_465(clk,rst,matrix2_A[17],matrix2_B[465],mul_res2[465]);
multi_7x41 multi_7x41_mod_466(clk,rst,matrix2_A[18],matrix2_B[466],mul_res2[466]);
multi_7x41 multi_7x41_mod_467(clk,rst,matrix2_A[19],matrix2_B[467],mul_res2[467]);
multi_7x41 multi_7x41_mod_468(clk,rst,matrix2_A[20],matrix2_B[468],mul_res2[468]);
multi_7x41 multi_7x41_mod_469(clk,rst,matrix2_A[21],matrix2_B[469],mul_res2[469]);
multi_7x41 multi_7x41_mod_470(clk,rst,matrix2_A[22],matrix2_B[470],mul_res2[470]);
multi_7x41 multi_7x41_mod_471(clk,rst,matrix2_A[23],matrix2_B[471],mul_res2[471]);
multi_7x41 multi_7x41_mod_472(clk,rst,matrix2_A[24],matrix2_B[472],mul_res2[472]);
multi_7x41 multi_7x41_mod_473(clk,rst,matrix2_A[25],matrix2_B[473],mul_res2[473]);
multi_7x41 multi_7x41_mod_474(clk,rst,matrix2_A[26],matrix2_B[474],mul_res2[474]);
multi_7x41 multi_7x41_mod_475(clk,rst,matrix2_A[27],matrix2_B[475],mul_res2[475]);
multi_7x41 multi_7x41_mod_476(clk,rst,matrix2_A[28],matrix2_B[476],mul_res2[476]);
multi_7x41 multi_7x41_mod_477(clk,rst,matrix2_A[29],matrix2_B[477],mul_res2[477]);
multi_7x41 multi_7x41_mod_478(clk,rst,matrix2_A[30],matrix2_B[478],mul_res2[478]);
multi_7x41 multi_7x41_mod_479(clk,rst,matrix2_A[31],matrix2_B[479],mul_res2[479]);
multi_7x41 multi_7x41_mod_480(clk,rst,matrix2_A[32],matrix2_B[480],mul_res2[480]);
multi_7x41 multi_7x41_mod_481(clk,rst,matrix2_A[33],matrix2_B[481],mul_res2[481]);
multi_7x41 multi_7x41_mod_482(clk,rst,matrix2_A[34],matrix2_B[482],mul_res2[482]);
multi_7x41 multi_7x41_mod_483(clk,rst,matrix2_A[35],matrix2_B[483],mul_res2[483]);
multi_7x41 multi_7x41_mod_484(clk,rst,matrix2_A[36],matrix2_B[484],mul_res2[484]);
multi_7x41 multi_7x41_mod_485(clk,rst,matrix2_A[37],matrix2_B[485],mul_res2[485]);
multi_7x41 multi_7x41_mod_486(clk,rst,matrix2_A[38],matrix2_B[486],mul_res2[486]);
multi_7x41 multi_7x41_mod_487(clk,rst,matrix2_A[39],matrix2_B[487],mul_res2[487]);
multi_7x41 multi_7x41_mod_488(clk,rst,matrix2_A[40],matrix2_B[488],mul_res2[488]);
multi_7x41 multi_7x41_mod_489(clk,rst,matrix2_A[41],matrix2_B[489],mul_res2[489]);
multi_7x41 multi_7x41_mod_490(clk,rst,matrix2_A[42],matrix2_B[490],mul_res2[490]);
multi_7x41 multi_7x41_mod_491(clk,rst,matrix2_A[43],matrix2_B[491],mul_res2[491]);
multi_7x41 multi_7x41_mod_492(clk,rst,matrix2_A[44],matrix2_B[492],mul_res2[492]);
multi_7x41 multi_7x41_mod_493(clk,rst,matrix2_A[45],matrix2_B[493],mul_res2[493]);
multi_7x41 multi_7x41_mod_494(clk,rst,matrix2_A[46],matrix2_B[494],mul_res2[494]);
multi_7x41 multi_7x41_mod_495(clk,rst,matrix2_A[47],matrix2_B[495],mul_res2[495]);
multi_7x41 multi_7x41_mod_496(clk,rst,matrix2_A[48],matrix2_B[496],mul_res2[496]);
multi_7x41 multi_7x41_mod_497(clk,rst,matrix2_A[49],matrix2_B[497],mul_res2[497]);
multi_7x41 multi_7x41_mod_498(clk,rst,matrix2_A[50],matrix2_B[498],mul_res2[498]);
multi_7x41 multi_7x41_mod_499(clk,rst,matrix2_A[51],matrix2_B[499],mul_res2[499]);
multi_7x41 multi_7x41_mod_500(clk,rst,matrix2_A[52],matrix2_B[500],mul_res2[500]);
multi_7x41 multi_7x41_mod_501(clk,rst,matrix2_A[53],matrix2_B[501],mul_res2[501]);
multi_7x41 multi_7x41_mod_502(clk,rst,matrix2_A[54],matrix2_B[502],mul_res2[502]);
multi_7x41 multi_7x41_mod_503(clk,rst,matrix2_A[55],matrix2_B[503],mul_res2[503]);
multi_7x41 multi_7x41_mod_504(clk,rst,matrix2_A[56],matrix2_B[504],mul_res2[504]);
multi_7x41 multi_7x41_mod_505(clk,rst,matrix2_A[57],matrix2_B[505],mul_res2[505]);
multi_7x41 multi_7x41_mod_506(clk,rst,matrix2_A[58],matrix2_B[506],mul_res2[506]);
multi_7x41 multi_7x41_mod_507(clk,rst,matrix2_A[59],matrix2_B[507],mul_res2[507]);
multi_7x41 multi_7x41_mod_508(clk,rst,matrix2_A[60],matrix2_B[508],mul_res2[508]);
multi_7x41 multi_7x41_mod_509(clk,rst,matrix2_A[61],matrix2_B[509],mul_res2[509]);
multi_7x41 multi_7x41_mod_510(clk,rst,matrix2_A[62],matrix2_B[510],mul_res2[510]);
multi_7x41 multi_7x41_mod_511(clk,rst,matrix2_A[63],matrix2_B[511],mul_res2[511]);
multi_7x41 multi_7x41_mod_512(clk,rst,matrix2_A[0],matrix2_B[512],mul_res2[512]);
multi_7x41 multi_7x41_mod_513(clk,rst,matrix2_A[1],matrix2_B[513],mul_res2[513]);
multi_7x41 multi_7x41_mod_514(clk,rst,matrix2_A[2],matrix2_B[514],mul_res2[514]);
multi_7x41 multi_7x41_mod_515(clk,rst,matrix2_A[3],matrix2_B[515],mul_res2[515]);
multi_7x41 multi_7x41_mod_516(clk,rst,matrix2_A[4],matrix2_B[516],mul_res2[516]);
multi_7x41 multi_7x41_mod_517(clk,rst,matrix2_A[5],matrix2_B[517],mul_res2[517]);
multi_7x41 multi_7x41_mod_518(clk,rst,matrix2_A[6],matrix2_B[518],mul_res2[518]);
multi_7x41 multi_7x41_mod_519(clk,rst,matrix2_A[7],matrix2_B[519],mul_res2[519]);
multi_7x41 multi_7x41_mod_520(clk,rst,matrix2_A[8],matrix2_B[520],mul_res2[520]);
multi_7x41 multi_7x41_mod_521(clk,rst,matrix2_A[9],matrix2_B[521],mul_res2[521]);
multi_7x41 multi_7x41_mod_522(clk,rst,matrix2_A[10],matrix2_B[522],mul_res2[522]);
multi_7x41 multi_7x41_mod_523(clk,rst,matrix2_A[11],matrix2_B[523],mul_res2[523]);
multi_7x41 multi_7x41_mod_524(clk,rst,matrix2_A[12],matrix2_B[524],mul_res2[524]);
multi_7x41 multi_7x41_mod_525(clk,rst,matrix2_A[13],matrix2_B[525],mul_res2[525]);
multi_7x41 multi_7x41_mod_526(clk,rst,matrix2_A[14],matrix2_B[526],mul_res2[526]);
multi_7x41 multi_7x41_mod_527(clk,rst,matrix2_A[15],matrix2_B[527],mul_res2[527]);
multi_7x41 multi_7x41_mod_528(clk,rst,matrix2_A[16],matrix2_B[528],mul_res2[528]);
multi_7x41 multi_7x41_mod_529(clk,rst,matrix2_A[17],matrix2_B[529],mul_res2[529]);
multi_7x41 multi_7x41_mod_530(clk,rst,matrix2_A[18],matrix2_B[530],mul_res2[530]);
multi_7x41 multi_7x41_mod_531(clk,rst,matrix2_A[19],matrix2_B[531],mul_res2[531]);
multi_7x41 multi_7x41_mod_532(clk,rst,matrix2_A[20],matrix2_B[532],mul_res2[532]);
multi_7x41 multi_7x41_mod_533(clk,rst,matrix2_A[21],matrix2_B[533],mul_res2[533]);
multi_7x41 multi_7x41_mod_534(clk,rst,matrix2_A[22],matrix2_B[534],mul_res2[534]);
multi_7x41 multi_7x41_mod_535(clk,rst,matrix2_A[23],matrix2_B[535],mul_res2[535]);
multi_7x41 multi_7x41_mod_536(clk,rst,matrix2_A[24],matrix2_B[536],mul_res2[536]);
multi_7x41 multi_7x41_mod_537(clk,rst,matrix2_A[25],matrix2_B[537],mul_res2[537]);
multi_7x41 multi_7x41_mod_538(clk,rst,matrix2_A[26],matrix2_B[538],mul_res2[538]);
multi_7x41 multi_7x41_mod_539(clk,rst,matrix2_A[27],matrix2_B[539],mul_res2[539]);
multi_7x41 multi_7x41_mod_540(clk,rst,matrix2_A[28],matrix2_B[540],mul_res2[540]);
multi_7x41 multi_7x41_mod_541(clk,rst,matrix2_A[29],matrix2_B[541],mul_res2[541]);
multi_7x41 multi_7x41_mod_542(clk,rst,matrix2_A[30],matrix2_B[542],mul_res2[542]);
multi_7x41 multi_7x41_mod_543(clk,rst,matrix2_A[31],matrix2_B[543],mul_res2[543]);
multi_7x41 multi_7x41_mod_544(clk,rst,matrix2_A[32],matrix2_B[544],mul_res2[544]);
multi_7x41 multi_7x41_mod_545(clk,rst,matrix2_A[33],matrix2_B[545],mul_res2[545]);
multi_7x41 multi_7x41_mod_546(clk,rst,matrix2_A[34],matrix2_B[546],mul_res2[546]);
multi_7x41 multi_7x41_mod_547(clk,rst,matrix2_A[35],matrix2_B[547],mul_res2[547]);
multi_7x41 multi_7x41_mod_548(clk,rst,matrix2_A[36],matrix2_B[548],mul_res2[548]);
multi_7x41 multi_7x41_mod_549(clk,rst,matrix2_A[37],matrix2_B[549],mul_res2[549]);
multi_7x41 multi_7x41_mod_550(clk,rst,matrix2_A[38],matrix2_B[550],mul_res2[550]);
multi_7x41 multi_7x41_mod_551(clk,rst,matrix2_A[39],matrix2_B[551],mul_res2[551]);
multi_7x41 multi_7x41_mod_552(clk,rst,matrix2_A[40],matrix2_B[552],mul_res2[552]);
multi_7x41 multi_7x41_mod_553(clk,rst,matrix2_A[41],matrix2_B[553],mul_res2[553]);
multi_7x41 multi_7x41_mod_554(clk,rst,matrix2_A[42],matrix2_B[554],mul_res2[554]);
multi_7x41 multi_7x41_mod_555(clk,rst,matrix2_A[43],matrix2_B[555],mul_res2[555]);
multi_7x41 multi_7x41_mod_556(clk,rst,matrix2_A[44],matrix2_B[556],mul_res2[556]);
multi_7x41 multi_7x41_mod_557(clk,rst,matrix2_A[45],matrix2_B[557],mul_res2[557]);
multi_7x41 multi_7x41_mod_558(clk,rst,matrix2_A[46],matrix2_B[558],mul_res2[558]);
multi_7x41 multi_7x41_mod_559(clk,rst,matrix2_A[47],matrix2_B[559],mul_res2[559]);
multi_7x41 multi_7x41_mod_560(clk,rst,matrix2_A[48],matrix2_B[560],mul_res2[560]);
multi_7x41 multi_7x41_mod_561(clk,rst,matrix2_A[49],matrix2_B[561],mul_res2[561]);
multi_7x41 multi_7x41_mod_562(clk,rst,matrix2_A[50],matrix2_B[562],mul_res2[562]);
multi_7x41 multi_7x41_mod_563(clk,rst,matrix2_A[51],matrix2_B[563],mul_res2[563]);
multi_7x41 multi_7x41_mod_564(clk,rst,matrix2_A[52],matrix2_B[564],mul_res2[564]);
multi_7x41 multi_7x41_mod_565(clk,rst,matrix2_A[53],matrix2_B[565],mul_res2[565]);
multi_7x41 multi_7x41_mod_566(clk,rst,matrix2_A[54],matrix2_B[566],mul_res2[566]);
multi_7x41 multi_7x41_mod_567(clk,rst,matrix2_A[55],matrix2_B[567],mul_res2[567]);
multi_7x41 multi_7x41_mod_568(clk,rst,matrix2_A[56],matrix2_B[568],mul_res2[568]);
multi_7x41 multi_7x41_mod_569(clk,rst,matrix2_A[57],matrix2_B[569],mul_res2[569]);
multi_7x41 multi_7x41_mod_570(clk,rst,matrix2_A[58],matrix2_B[570],mul_res2[570]);
multi_7x41 multi_7x41_mod_571(clk,rst,matrix2_A[59],matrix2_B[571],mul_res2[571]);
multi_7x41 multi_7x41_mod_572(clk,rst,matrix2_A[60],matrix2_B[572],mul_res2[572]);
multi_7x41 multi_7x41_mod_573(clk,rst,matrix2_A[61],matrix2_B[573],mul_res2[573]);
multi_7x41 multi_7x41_mod_574(clk,rst,matrix2_A[62],matrix2_B[574],mul_res2[574]);
multi_7x41 multi_7x41_mod_575(clk,rst,matrix2_A[63],matrix2_B[575],mul_res2[575]);
multi_7x41 multi_7x41_mod_576(clk,rst,matrix2_A[0],matrix2_B[576],mul_res2[576]);
multi_7x41 multi_7x41_mod_577(clk,rst,matrix2_A[1],matrix2_B[577],mul_res2[577]);
multi_7x41 multi_7x41_mod_578(clk,rst,matrix2_A[2],matrix2_B[578],mul_res2[578]);
multi_7x41 multi_7x41_mod_579(clk,rst,matrix2_A[3],matrix2_B[579],mul_res2[579]);
multi_7x41 multi_7x41_mod_580(clk,rst,matrix2_A[4],matrix2_B[580],mul_res2[580]);
multi_7x41 multi_7x41_mod_581(clk,rst,matrix2_A[5],matrix2_B[581],mul_res2[581]);
multi_7x41 multi_7x41_mod_582(clk,rst,matrix2_A[6],matrix2_B[582],mul_res2[582]);
multi_7x41 multi_7x41_mod_583(clk,rst,matrix2_A[7],matrix2_B[583],mul_res2[583]);
multi_7x41 multi_7x41_mod_584(clk,rst,matrix2_A[8],matrix2_B[584],mul_res2[584]);
multi_7x41 multi_7x41_mod_585(clk,rst,matrix2_A[9],matrix2_B[585],mul_res2[585]);
multi_7x41 multi_7x41_mod_586(clk,rst,matrix2_A[10],matrix2_B[586],mul_res2[586]);
multi_7x41 multi_7x41_mod_587(clk,rst,matrix2_A[11],matrix2_B[587],mul_res2[587]);
multi_7x41 multi_7x41_mod_588(clk,rst,matrix2_A[12],matrix2_B[588],mul_res2[588]);
multi_7x41 multi_7x41_mod_589(clk,rst,matrix2_A[13],matrix2_B[589],mul_res2[589]);
multi_7x41 multi_7x41_mod_590(clk,rst,matrix2_A[14],matrix2_B[590],mul_res2[590]);
multi_7x41 multi_7x41_mod_591(clk,rst,matrix2_A[15],matrix2_B[591],mul_res2[591]);
multi_7x41 multi_7x41_mod_592(clk,rst,matrix2_A[16],matrix2_B[592],mul_res2[592]);
multi_7x41 multi_7x41_mod_593(clk,rst,matrix2_A[17],matrix2_B[593],mul_res2[593]);
multi_7x41 multi_7x41_mod_594(clk,rst,matrix2_A[18],matrix2_B[594],mul_res2[594]);
multi_7x41 multi_7x41_mod_595(clk,rst,matrix2_A[19],matrix2_B[595],mul_res2[595]);
multi_7x41 multi_7x41_mod_596(clk,rst,matrix2_A[20],matrix2_B[596],mul_res2[596]);
multi_7x41 multi_7x41_mod_597(clk,rst,matrix2_A[21],matrix2_B[597],mul_res2[597]);
multi_7x41 multi_7x41_mod_598(clk,rst,matrix2_A[22],matrix2_B[598],mul_res2[598]);
multi_7x41 multi_7x41_mod_599(clk,rst,matrix2_A[23],matrix2_B[599],mul_res2[599]);
multi_7x41 multi_7x41_mod_600(clk,rst,matrix2_A[24],matrix2_B[600],mul_res2[600]);
multi_7x41 multi_7x41_mod_601(clk,rst,matrix2_A[25],matrix2_B[601],mul_res2[601]);
multi_7x41 multi_7x41_mod_602(clk,rst,matrix2_A[26],matrix2_B[602],mul_res2[602]);
multi_7x41 multi_7x41_mod_603(clk,rst,matrix2_A[27],matrix2_B[603],mul_res2[603]);
multi_7x41 multi_7x41_mod_604(clk,rst,matrix2_A[28],matrix2_B[604],mul_res2[604]);
multi_7x41 multi_7x41_mod_605(clk,rst,matrix2_A[29],matrix2_B[605],mul_res2[605]);
multi_7x41 multi_7x41_mod_606(clk,rst,matrix2_A[30],matrix2_B[606],mul_res2[606]);
multi_7x41 multi_7x41_mod_607(clk,rst,matrix2_A[31],matrix2_B[607],mul_res2[607]);
multi_7x41 multi_7x41_mod_608(clk,rst,matrix2_A[32],matrix2_B[608],mul_res2[608]);
multi_7x41 multi_7x41_mod_609(clk,rst,matrix2_A[33],matrix2_B[609],mul_res2[609]);
multi_7x41 multi_7x41_mod_610(clk,rst,matrix2_A[34],matrix2_B[610],mul_res2[610]);
multi_7x41 multi_7x41_mod_611(clk,rst,matrix2_A[35],matrix2_B[611],mul_res2[611]);
multi_7x41 multi_7x41_mod_612(clk,rst,matrix2_A[36],matrix2_B[612],mul_res2[612]);
multi_7x41 multi_7x41_mod_613(clk,rst,matrix2_A[37],matrix2_B[613],mul_res2[613]);
multi_7x41 multi_7x41_mod_614(clk,rst,matrix2_A[38],matrix2_B[614],mul_res2[614]);
multi_7x41 multi_7x41_mod_615(clk,rst,matrix2_A[39],matrix2_B[615],mul_res2[615]);
multi_7x41 multi_7x41_mod_616(clk,rst,matrix2_A[40],matrix2_B[616],mul_res2[616]);
multi_7x41 multi_7x41_mod_617(clk,rst,matrix2_A[41],matrix2_B[617],mul_res2[617]);
multi_7x41 multi_7x41_mod_618(clk,rst,matrix2_A[42],matrix2_B[618],mul_res2[618]);
multi_7x41 multi_7x41_mod_619(clk,rst,matrix2_A[43],matrix2_B[619],mul_res2[619]);
multi_7x41 multi_7x41_mod_620(clk,rst,matrix2_A[44],matrix2_B[620],mul_res2[620]);
multi_7x41 multi_7x41_mod_621(clk,rst,matrix2_A[45],matrix2_B[621],mul_res2[621]);
multi_7x41 multi_7x41_mod_622(clk,rst,matrix2_A[46],matrix2_B[622],mul_res2[622]);
multi_7x41 multi_7x41_mod_623(clk,rst,matrix2_A[47],matrix2_B[623],mul_res2[623]);
multi_7x41 multi_7x41_mod_624(clk,rst,matrix2_A[48],matrix2_B[624],mul_res2[624]);
multi_7x41 multi_7x41_mod_625(clk,rst,matrix2_A[49],matrix2_B[625],mul_res2[625]);
multi_7x41 multi_7x41_mod_626(clk,rst,matrix2_A[50],matrix2_B[626],mul_res2[626]);
multi_7x41 multi_7x41_mod_627(clk,rst,matrix2_A[51],matrix2_B[627],mul_res2[627]);
multi_7x41 multi_7x41_mod_628(clk,rst,matrix2_A[52],matrix2_B[628],mul_res2[628]);
multi_7x41 multi_7x41_mod_629(clk,rst,matrix2_A[53],matrix2_B[629],mul_res2[629]);
multi_7x41 multi_7x41_mod_630(clk,rst,matrix2_A[54],matrix2_B[630],mul_res2[630]);
multi_7x41 multi_7x41_mod_631(clk,rst,matrix2_A[55],matrix2_B[631],mul_res2[631]);
multi_7x41 multi_7x41_mod_632(clk,rst,matrix2_A[56],matrix2_B[632],mul_res2[632]);
multi_7x41 multi_7x41_mod_633(clk,rst,matrix2_A[57],matrix2_B[633],mul_res2[633]);
multi_7x41 multi_7x41_mod_634(clk,rst,matrix2_A[58],matrix2_B[634],mul_res2[634]);
multi_7x41 multi_7x41_mod_635(clk,rst,matrix2_A[59],matrix2_B[635],mul_res2[635]);
multi_7x41 multi_7x41_mod_636(clk,rst,matrix2_A[60],matrix2_B[636],mul_res2[636]);
multi_7x41 multi_7x41_mod_637(clk,rst,matrix2_A[61],matrix2_B[637],mul_res2[637]);
multi_7x41 multi_7x41_mod_638(clk,rst,matrix2_A[62],matrix2_B[638],mul_res2[638]);
multi_7x41 multi_7x41_mod_639(clk,rst,matrix2_A[63],matrix2_B[639],mul_res2[639]);


/*

#include <stdio.h>
   
   int main() {
       // Write C code here
       int i,j;
       int k = 0;
       int z = 0;
      
        for (j = 0; j<10;j++) { // columns
          for(i =0; i<64; i++){    //64-1 rows

            z = ((10 * i) - 1 + j) < 0 ? 0 : ((10 * i)  + j); // 10 is width of matrix
            
printf("multi_7x41 multi_7x41_mod_%d(clk,rst,matrix2_A[%d],matrix2_B[%d],mul_res2[%d]);\n",k,i,k,k);
k = k+1;



  }
}
       return 0;
   }



*/

adder_64in adder_64in_mod_0(clk,rst,mul_res2[0], mul_res2[1], mul_res2[2], mul_res2[3], mul_res2[4], mul_res2[5], mul_res2[6], mul_res2[7], mul_res2[8], mul_res2[9], mul_res2[10], mul_res2[11], mul_res2[12], mul_res2[13], mul_res2[14], mul_res2[15], mul_res2[16], mul_res2[17], mul_res2[18], mul_res2[19], mul_res2[20], mul_res2[21], mul_res2[22], mul_res2[23], mul_res2[24], mul_res2[25], mul_res2[26], mul_res2[27], mul_res2[28], mul_res2[29], mul_res2[30], mul_res2[31], mul_res2[32], mul_res2[33], mul_res2[34], mul_res2[35], mul_res2[36], mul_res2[37], mul_res2[38], mul_res2[39], mul_res2[40], mul_res2[41], mul_res2[42], mul_res2[43], mul_res2[44], mul_res2[45], mul_res2[46], mul_res2[47], mul_res2[48], mul_res2[49], mul_res2[50], mul_res2[51], mul_res2[52], mul_res2[53], mul_res2[54], mul_res2[55], mul_res2[56], mul_res2[57], mul_res2[58], mul_res2[59], mul_res2[60], mul_res2[61], mul_res2[62], mul_res2[63],result_fc2[0]);


adder_64in adder_64in_mod_1(clk,rst,mul_res2[64], mul_res2[65], mul_res2[66], mul_res2[67], mul_res2[68], mul_res2[69], mul_res2[70], mul_res2[71], mul_res2[72], mul_res2[73], mul_res2[74], mul_res2[75], mul_res2[76], mul_res2[77], mul_res2[78], mul_res2[79], mul_res2[80], mul_res2[81], mul_res2[82], mul_res2[83], mul_res2[84], mul_res2[85], mul_res2[86], mul_res2[87], mul_res2[88], mul_res2[89], mul_res2[90], mul_res2[91], mul_res2[92], mul_res2[93], mul_res2[94], mul_res2[95], mul_res2[96], mul_res2[97], mul_res2[98], mul_res2[99], mul_res2[100], mul_res2[101], mul_res2[102], mul_res2[103], mul_res2[104], mul_res2[105], mul_res2[106], mul_res2[107], mul_res2[108], mul_res2[109], mul_res2[110], mul_res2[111], mul_res2[112], mul_res2[113], mul_res2[114], mul_res2[115], mul_res2[116], mul_res2[117], mul_res2[118], mul_res2[119], mul_res2[120], mul_res2[121], mul_res2[122], mul_res2[123], mul_res2[124], mul_res2[125], mul_res2[126], mul_res2[127],result_fc2[1]);


adder_64in adder_64in_mod_2(clk,rst,mul_res2[128], mul_res2[129], mul_res2[130], mul_res2[131], mul_res2[132], mul_res2[133], mul_res2[134], mul_res2[135], mul_res2[136], mul_res2[137], mul_res2[138], mul_res2[139], mul_res2[140], mul_res2[141], mul_res2[142], mul_res2[143], mul_res2[144], mul_res2[145], mul_res2[146], mul_res2[147], mul_res2[148], mul_res2[149], mul_res2[150], mul_res2[151], mul_res2[152], mul_res2[153], mul_res2[154], mul_res2[155], mul_res2[156], mul_res2[157], mul_res2[158], mul_res2[159], mul_res2[160], mul_res2[161], mul_res2[162], mul_res2[163], mul_res2[164], mul_res2[165], mul_res2[166], mul_res2[167], mul_res2[168], mul_res2[169], mul_res2[170], mul_res2[171], mul_res2[172], mul_res2[173], mul_res2[174], mul_res2[175], mul_res2[176], mul_res2[177], 
mul_res2[178], mul_res2[179], mul_res2[180], mul_res2[181], mul_res2[182], mul_res2[183], mul_res2[184], mul_res2[185], mul_res2[186], mul_res2[187], mul_res2[188], mul_res2[189], mul_res2[190], mul_res2[191],result_fc2[2]);


adder_64in adder_64in_mod_3(clk,rst,mul_res2[192], mul_res2[193], mul_res2[194], mul_res2[195], mul_res2[196], mul_res2[197], mul_res2[198], mul_res2[199], mul_res2[200], mul_res2[201], mul_res2[202], mul_res2[203], mul_res2[204], mul_res2[205], mul_res2[206], mul_res2[207], mul_res2[208], mul_res2[209], mul_res2[210], mul_res2[211], mul_res2[212], mul_res2[213], mul_res2[214], mul_res2[215], mul_res2[216], mul_res2[217], mul_res2[218], mul_res2[219], mul_res2[220], mul_res2[221], mul_res2[222], mul_res2[223], mul_res2[224], mul_res2[225], mul_res2[226], mul_res2[227], mul_res2[228], mul_res2[229], mul_res2[230], mul_res2[231], mul_res2[232], mul_res2[233], mul_res2[234], mul_res2[235], mul_res2[236], mul_res2[237], mul_res2[238], mul_res2[239], mul_res2[240], mul_res2[241], 
mul_res2[242], mul_res2[243], mul_res2[244], mul_res2[245], mul_res2[246], mul_res2[247], mul_res2[248], mul_res2[249], mul_res2[250], mul_res2[251], mul_res2[252], mul_res2[253], mul_res2[254], mul_res2[255],result_fc2[3]);


adder_64in adder_64in_mod_4(clk,rst,mul_res2[256], mul_res2[257], mul_res2[258], mul_res2[259], mul_res2[260], mul_res2[261], mul_res2[262], mul_res2[263], mul_res2[264], mul_res2[265], mul_res2[266], mul_res2[267], mul_res2[268], mul_res2[269], mul_res2[270], mul_res2[271], mul_res2[272], mul_res2[273], mul_res2[274], mul_res2[275], mul_res2[276], mul_res2[277], mul_res2[278], mul_res2[279], mul_res2[280], mul_res2[281], mul_res2[282], mul_res2[283], mul_res2[284], mul_res2[285], mul_res2[286], mul_res2[287], mul_res2[288], mul_res2[289], mul_res2[290], mul_res2[291], mul_res2[292], mul_res2[293], mul_res2[294], mul_res2[295], mul_res2[296], mul_res2[297], mul_res2[298], mul_res2[299], mul_res2[300], mul_res2[301], mul_res2[302], mul_res2[303], mul_res2[304], mul_res2[305], 
mul_res2[306], mul_res2[307], mul_res2[308], mul_res2[309], mul_res2[310], mul_res2[311], mul_res2[312], mul_res2[313], mul_res2[314], mul_res2[315], mul_res2[316], mul_res2[317], mul_res2[318], mul_res2[319],result_fc2[4]);


adder_64in adder_64in_mod_5(clk,rst,mul_res2[320], mul_res2[321], mul_res2[322], mul_res2[323], mul_res2[324], mul_res2[325], mul_res2[326], mul_res2[327], mul_res2[328], mul_res2[329], mul_res2[330], mul_res2[331], mul_res2[332], mul_res2[333], mul_res2[334], mul_res2[335], mul_res2[336], mul_res2[337], mul_res2[338], mul_res2[339], mul_res2[340], mul_res2[341], mul_res2[342], mul_res2[343], mul_res2[344], mul_res2[345], mul_res2[346], mul_res2[347], mul_res2[348], mul_res2[349], mul_res2[350], mul_res2[351], mul_res2[352], mul_res2[353], mul_res2[354], mul_res2[355], mul_res2[356], mul_res2[357], mul_res2[358], mul_res2[359], mul_res2[360], mul_res2[361], mul_res2[362], mul_res2[363], mul_res2[364], mul_res2[365], mul_res2[366], mul_res2[367], mul_res2[368], mul_res2[369], 
mul_res2[370], mul_res2[371], mul_res2[372], mul_res2[373], mul_res2[374], mul_res2[375], mul_res2[376], mul_res2[377], mul_res2[378], mul_res2[379], mul_res2[380], mul_res2[381], mul_res2[382], mul_res2[383],result_fc2[5]);


adder_64in adder_64in_mod_6(clk,rst,mul_res2[384], mul_res2[385], mul_res2[386], mul_res2[387], mul_res2[388], mul_res2[389], mul_res2[390], mul_res2[391], mul_res2[392], mul_res2[393], mul_res2[394], mul_res2[395], mul_res2[396], mul_res2[397], mul_res2[398], mul_res2[399], mul_res2[400], mul_res2[401], mul_res2[402], mul_res2[403], mul_res2[404], mul_res2[405], mul_res2[406], mul_res2[407], mul_res2[408], mul_res2[409], mul_res2[410], mul_res2[411], mul_res2[412], mul_res2[413], mul_res2[414], mul_res2[415], mul_res2[416], mul_res2[417], mul_res2[418], mul_res2[419], mul_res2[420], mul_res2[421], mul_res2[422], mul_res2[423], mul_res2[424], mul_res2[425], mul_res2[426], mul_res2[427], mul_res2[428], mul_res2[429], mul_res2[430], mul_res2[431], mul_res2[432], mul_res2[433], 
mul_res2[434], mul_res2[435], mul_res2[436], mul_res2[437], mul_res2[438], mul_res2[439], mul_res2[440], mul_res2[441], mul_res2[442], mul_res2[443], mul_res2[444], mul_res2[445], mul_res2[446], mul_res2[447],result_fc2[6]);


adder_64in adder_64in_mod_7(clk,rst,mul_res2[448], mul_res2[449], mul_res2[450], mul_res2[451], mul_res2[452], mul_res2[453], mul_res2[454], mul_res2[455], mul_res2[456], mul_res2[457], mul_res2[458], mul_res2[459], mul_res2[460], mul_res2[461], mul_res2[462], mul_res2[463], mul_res2[464], mul_res2[465], mul_res2[466], mul_res2[467], mul_res2[468], mul_res2[469], mul_res2[470], mul_res2[471], mul_res2[472], mul_res2[473], mul_res2[474], mul_res2[475], mul_res2[476], mul_res2[477], mul_res2[478], mul_res2[479], mul_res2[480], mul_res2[481], mul_res2[482], mul_res2[483], mul_res2[484], mul_res2[485], mul_res2[486], mul_res2[487], mul_res2[488], mul_res2[489], mul_res2[490], mul_res2[491], mul_res2[492], mul_res2[493], mul_res2[494], mul_res2[495], mul_res2[496], mul_res2[497], 
mul_res2[498], mul_res2[499], mul_res2[500], mul_res2[501], mul_res2[502], mul_res2[503], mul_res2[504], mul_res2[505], mul_res2[506], mul_res2[507], mul_res2[508], mul_res2[509], mul_res2[510], mul_res2[511],result_fc2[7]);


adder_64in adder_64in_mod_8(clk,rst,mul_res2[512], mul_res2[513], mul_res2[514], mul_res2[515], mul_res2[516], mul_res2[517], mul_res2[518], mul_res2[519], mul_res2[520], mul_res2[521], mul_res2[522], mul_res2[523], mul_res2[524], mul_res2[525], mul_res2[526], mul_res2[527], mul_res2[528], mul_res2[529], mul_res2[530], mul_res2[531], mul_res2[532], mul_res2[533], mul_res2[534], mul_res2[535], mul_res2[536], mul_res2[537], mul_res2[538], mul_res2[539], mul_res2[540], mul_res2[541], mul_res2[542], mul_res2[543], mul_res2[544], mul_res2[545], mul_res2[546], mul_res2[547], mul_res2[548], mul_res2[549], mul_res2[550], mul_res2[551], mul_res2[552], mul_res2[553], mul_res2[554], mul_res2[555], mul_res2[556], mul_res2[557], mul_res2[558], mul_res2[559], mul_res2[560], mul_res2[561], 
mul_res2[562], mul_res2[563], mul_res2[564], mul_res2[565], mul_res2[566], mul_res2[567], mul_res2[568], mul_res2[569], mul_res2[570], mul_res2[571], mul_res2[572], mul_res2[573], mul_res2[574], mul_res2[575],result_fc2[8]);


adder_64in adder_64in_mod_9(clk,rst,mul_res2[576], mul_res2[577], mul_res2[578], mul_res2[579], mul_res2[580], mul_res2[581], mul_res2[582], mul_res2[583], mul_res2[584], mul_res2[585], mul_res2[586], mul_res2[587], mul_res2[588], mul_res2[589], mul_res2[590], mul_res2[591], mul_res2[592], mul_res2[593], mul_res2[594], mul_res2[595], mul_res2[596], mul_res2[597], mul_res2[598], mul_res2[599], mul_res2[600], mul_res2[601], mul_res2[602], mul_res2[603], mul_res2[604], mul_res2[605], mul_res2[606], mul_res2[607], mul_res2[608], mul_res2[609], mul_res2[610], mul_res2[611], mul_res2[612], mul_res2[613], mul_res2[614], mul_res2[615], mul_res2[616], mul_res2[617], mul_res2[618], mul_res2[619], mul_res2[620], mul_res2[621], mul_res2[622], mul_res2[623], mul_res2[624], mul_res2[625], 
mul_res2[626], mul_res2[627], mul_res2[628], mul_res2[629], mul_res2[630], mul_res2[631], mul_res2[632], mul_res2[633], mul_res2[634], mul_res2[635], mul_res2[636], mul_res2[637], mul_res2[638], mul_res2[639],result_fc2[9]);



endmodule
