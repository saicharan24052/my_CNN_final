

// convert it to kernel_1_re[4][9]
  reg  signed [7:0] kernel_1_re [4][9] = '{
  '{68, 56, 32, 66, 78, 67, 53, 65, 77},
  '{75, 65, 43, 63, 76, 61, 35, 56, 71},
  '{74, 62, 39, 66, 76, 65, 48, 62, 73},
  '{69, 64, 47, 63, 80, 73, 40, 56, 64}
};


//////////////////////////////
/*
 real kernel_1_re[4][3][3] = '{
  '{
    '{
      '{39, 37, 38},
      '{47, 47, 44},
      '{42, 43, 36} 
    } 
  },
  '{
    '{
      '{40, 41, 33},
      '{48, 54, 46},
      '{39, 40, 41} 
    } 
  },
  '{
    '{
      '{31, 37, 38},
      '{45, 48, 44},
      '{40, 45, 40} 
    } 
  },
  '{
    '{
      '{37, 43, 36},
      '{41, 47, 47},
      '{42, 43, 41} 
    } 
  } 
};
*/
/*
 real kernel_2_re[8][3][3] = '{
  '{
    '{
      '{-8, -49, -59},
      '{40, 22, 15},
      '{29, 26, 35} 
    },
    '{
      '{-4, -44, -59},
      '{43, 22, 20},
      '{28, 29, 37} 
    },
    '{
      '{0, -43, -55},
      '{42, 20, 26},
      '{26, 26, 38} 
    },
    '{
      '{-4, -42, -59},
      '{35, 24, 24},
      '{27, 30, 42} 
    } 
  },
  '{
    '{
      '{36, 43, 50},
      '{-10, -2, -12},
      '{-59, -53, -43} 
    },
    '{
      '{37, 42, 52},
      '{-5, -4, -9},
      '{-58, -52, -46} 
    },
    '{
      '{40, 45, 44},
      '{-7, 1, -13},
      '{-55, -48, -33} 
    },
    '{
      '{33, 45, 49},
      '{-6, -1, -8},
      '{-61, -53, -48} 
    } 
  },
  '{
    '{
      '{29, 44, 33},
      '{-35, -6, 31},
      '{-27, -1, 35} 
    },
    '{
      '{26, 42, 42},
      '{-36, -8, 32},
      '{-25, -1, 33} 
    },
    '{
      '{29, 42, 36},
      '{-25, -3, 35},
      '{-26, 10, 41} 
    },
    '{
      '{30, 41, 36},
      '{-33, -4, 31},
      '{-25, -1, 36} 
    } 
  },
  '{
    '{
      '{-56, -7, 44},
      '{-61, 20, 37},
      '{-23, 27, 29} 
    },
    '{
      '{-60, -1, 48},
      '{-60, 26, 32},
      '{-29, 25, 23} 
    },
    '{
      '{-58, -4, 44},
      '{-61, 18, 33},
      '{-26, 30, 23} 
    },
    '{
      '{-62, -2, 48},
      '{-55, 24, 33},
      '{-25, 31, 24} 
    } 
  },
  '{
    '{
      '{23, 20, 18},
      '{20, 18, 7},
      '{19, 15, 20} 
    },
    '{
      '{20, 21, 28},
      '{13, 11, 10},
      '{21, 4, 18} 
    },
    '{
      '{26, 26, 19},
      '{15, 13, 8},
      '{16, 10, 14} 
    },
    '{
      '{21, 24, 19},
      '{13, 13, 8},
      '{16, 15, 14} 
    } 
  },
  '{
    '{
      '{22, 23, 24},
      '{18, 28, 42},
      '{-57, -54, -20} 
    },
    '{
      '{30, 23, 29},
      '{18, 28, 38},
      '{-57, -53, -16} 
    },
    '{
      '{27, 23, 29},
      '{22, 25, 44},
      '{-54, -55, -16} 
    },
    '{
      '{29, 24, 25},
      '{14, 27, 44},
      '{-57, -56, -11} 
    } 
  },
  '{
    '{
      '{-19, 15, 31},
      '{27, 24, 25},
      '{28, 17, 5} 
    },
    '{
      '{-18, 9, 34},
      '{26, 22, 22},
      '{27, 19, -1} 
    },
    '{
      '{-16, 20, 36},
      '{34, 26, 24},
      '{34, 20, -6} 
    },
    '{
      '{-14, 19, 36},
      '{29, 26, 21},
      '{27, 14, 0} 
    } 
  },
  '{
    '{
      '{10, 22, 23},
      '{16, 20, 12},
      '{24, 20, 25} 
    },
    '{
      '{8, 23, 27},
      '{18, 15, 20},
      '{22, 19, 22} 
    },
    '{
      '{16, 22, 20},
      '{21, 22, 9},
      '{20, 19, 17} 
    },
    '{
      '{16, 23, 28},
      '{19, 20, 13},
      '{20, 20, 24} 
    } 
  } 
};
*/
  reg  signed [7:0] kernel_2_re[32][9] ='{
  '{3, 27, 21, 31, 9, 5, 49, 12, 10},
  '{8, 29, 21, 33, 16, 3, 47, 8, 7},
  '{2, 34, 19, 33, 13, 0, 46, 7, 2},
  '{8, 34, 20, 33, 11, 4, 53, 8, 10},

  '{-6, 42, 42, -75, 24, 55, -118, -1, 62},
  '{-1, 46, 42, -78, 30, 63, -113, 10, 61},
  '{-5, 46, 52, -80, 27, 55, -115, -1, 61},
  '{-5, 40, 44, -78, 24, 56, -119, 2, 51},

  '{-63, 21, 48, -27, 53, 26, 61, 53, 13},
  '{-61, 21, 45, -27, 50, 30, 53, 53, 8},
  '{-61, 13, 51, -30, 57, 27, 59, 57, 14},
  '{-63, 17, 53, -38, 53, 33, 55, 56, 10},

  '{34, 29, -8, 3, 40, 37, -54, 0, 27},
  '{40, 33, -3, 11, 43, 38, -51, 6, 30},
  '{34, 32, -6, 6, 40, 37, -59, 2, 33},
  '{36, 29, -3, 8, 38, 30, -56, 6, 37},

  '{2, -89, -108, 75, 51, 28, 51, 57, 69},
  '{-4, -92, -104, 73, 45, 26, 50, 57, 73},
  '{4, -89, -110, 73, 47, 26, 46, 54, 67},
  '{-4, -92, -112, 72, 30, 14, 43, 57, 70},

  '{38, 36, 56, 32, 45, 52, -97, -93, -63},
  '{36, 26, 45, 41, 47, 62, -94, -90, -61},
  '{36, 39, 49, 40, 56, 54, -93, -94, -66},
  '{34, 36, 51, 45, 57, 63, -90, -97, -60},

  '{-17, 7, 38, 29, 24, 46, 38, 19, 39},
  '{-20, 5, 35, 23, 31, 39, 37, 20, 43},
  '{-30, 4, 35, 24, 30, 45, 36, 16, 42},
  '{-28, 2, 42, 21, 27, 42, 33, 19, 44},

  '{38, 40, -4, 3, 30, 7, -19, 45, 43},
  '{44, 49, -2, 14, 34, 3, -19, 46, 49},
  '{40, 44, 1, 6, 24, 0, -19, 43, 46},
  '{42, 45, 2, 5, 30, 2, -19, 41, 44}
};

 
 /*
// 7 bit without sign
reg  signed [7:0] fc1_weights_re[64][200] = '{
  '{4, 42, -2, -5, -1, -5, -23, -46, -39, -14, -8, 22, 47, 12, 21, -4, 39, 34, 17, -26, -37, 0, 14, 23, -5, -29, 4, -5, 7, -49, -25, -12, 37, -9, -71, 43, -9, 7, -34, 33, -23, -18, 25, -12, -11, -37, 15, 8, -4, 8, 11, -16, 0, -42, -13, -14, -13, -12, 61, 26, 6, 5, 17, -15, 20, 25, -20, -30, 40, -46, -9, 31, 16, 27, -1, -5, -34, 23, -28, -46, -30, 10, -38, -29, -34, -3, -40, -42, -8, 27, 15, 20, -4, -37, -9, -33, -6, -45, -57, 29, -8, 28, -11, 41, -24, 5, 8, 4, -27, 5, -20, 24, -35, -9, 49, 41, -22, 20, 26, -18, 14, 51, 27, 44, 19, -28, 19, 66, 49, 14, 36, -2, 53, 42, 8, -34, -16, 19, -37, 36, 4, -34, 1, 14, 14, 19, -3, -37, 28, 9, -19, 38, 0, 47, 9, 30, 33, 19, 1, 10, 11, -10, -7, -21, -7, 5, -4, -3, 8, -17, 18, 37, -32, -3, 0, 32, -1, 13, 54, 31, -38, -33, 33, -35, 36, 36, -17, -5, 13, 52, -15, 39, -22, 6, 36, 44, 2, -17, -9, 33},
  '{2, 32, 7, 51, 51, 25, 5, 25, 20, 7, 42, 38, -14, -36, -18, 12, -4, -24, -11, -7, -43, -50, -7, -35, -1, -14, -4, 29, -28, -31, -22, 4, 31, 11, -49, -6, -19, -17, -21, 4, -40, -18, 21, 28, 31, -29, 28, 26, 23, -17, -24, -11, 11, -16, -9, -8, 5, -11, 21, 14, 7, 11, 19, 35, -42, -4, -23, -23, -20, -46, 21, -11, 12, -32, 53, -7, -11, -23, -21, -24, 22, 18, -16, 13, 20, -12, -1, -33, 37, 41, -7, -6, -14, 0, -33, 13, -4, -5, 8, -18, 22, 24, -24, -12, 7, 15, 11, 26, -14, -9, -21, -10, 26, 14, 38, 45, 21, 36, -17, -24, -15, 28, -7, 19, 24, -8, -37, 6, 8, -42, 6, 34, -14, 36, 12, 26, 60, 31, 11, 29, 6, 47, -17, 37, 2, -23, 16, -32, -20, 17, -12, 31, 28, -6, 8, 33, 44, -5, 12, 18, -11, 2, -6, 41, 11, 51, 43, -25, 53, -29, -28, 21, -40, 4, 20, -10, 47, -14, 13, -20, 16, -17, 26, -8, 36, 3, 10, -40, 27, 16, 20, 16, 10, 8, -1, -30, -34, -48, 31, 10},
  '{-17, 20, -32, 10, 21, -12, 49, -4, 3, 18, 33, 7, -12, 22, 24, 30, 35, 3, 30, 32, 22, -3, 60, 31, -8, -3, 11, -38, 13, 52, 25, -21, 15, 4, 83, -37, -1, 43, 58, -23, 0, 20, 10, 4, -73, 33, -17, -22, -4, -6, 18, -6, 30, -7, -15, -18, -13, -1, -28, -32, 12, -27, -37, -18, 12, -17, -20, -25, 16, -7, 21, 9, -10, -23, -35, 18, -16, 13, -1, 0, -3, 5, 24, 3, -6, -19, 16, 7, -38, -51, -36, 9, 4, 35, 15, -15, 32, -7, 40, 23, 8, 11, -15, 0, -16, 36, -27, -18, 29, -18, 37, 49, -25, 19, -4, 1, -30, -20, -48, 29, 13, 16, -9, 3, 18, 16, 34, -22, 29, -10, 25, -40, -25, 35, 35, -16, -16, 40, 2, 16, -3, 47, 0, -22, -19, 19, -28, -14, -10, -8, 26, -37, -7, -4, 17, -21, -4, 17, 9, -3, -12, 34, 39, -34, 17, 11, -6, -23, -29, -12, 30, 13, 6, 5, -2, 11, 0, -10, -9, 19, -22, 12, 46, -26, -33, 21, 24, 28, -40, -21, -29, 3, -20, 5, 41, -36, -7, 27, -5, 25},
  '{-1, -9, -11, 25, 33, 5, 43, -5, 8, 21, 15, -21, 15, 50, 25, 5, 9, 36, 3, 4, -14, -29, -28, -19, -18, 28, -42, 14, 83, 82, -36, -25, 49, 45, 60, -27, 3, 46, 20, 46, 23, 9, 9, 22, -21, 20, 63, 0, 19, -9, 23, 24, -16, -10, 17, 21, -8, -7, -30, 4, 29, 24, 35, -21, -15, -3, 15, 30, 2, 43, 37, 2, 38, -19, 36, -6, -18, -9, 4, -7, 37, 21, 3, -33, -43, -17, 1, 23, -29, -23, -10, -38, 12, 31, 11, 26, -1, 19, -6, 31, 8, 17, -23, 7, -41, 43, -17, 37, 8, -16, 3, 32, -14, -16, -13, -35, -22, -14, 32, -34, -29, -8, 25, -17, 12, 4, -2, -51, -27, 21, -52, -45, -14, 2, 19, -15, 23, -16, -4, 20, 32, -5, -9, 1, 2, -32, 23, 28, 6, -40, -40, 14, 9, -1, -35, 22, 39, 24, -13, -35, 26, -36, -11, -2, 27, 10, -6, -15, -23, -44, 33, 1, 41, -5, -28, -22, -36, 16, 18, 3, 21, -18, 12, 42, 12, -12, 34, 47, 33, 23, -21, -2, -19, -18, -14, -21, 8, 53, -25, -15},
  '{39, -31, 17, 44, 11, -8, -15, -9, 52, 16, -37, -38, 32, 9, 31, 7, 40, 14, -38, 27, 72, 71, -7, -6, -47, 19, 19, 30, 29, 49, -36, -18, -1, -9, 11, -23, -8, 17, 6, 23, 36, 43, 16, -17, -57, 63, 22, -9, -15, -4, -30, 4, -37, -15, -1, 2, 7, 2, -23, 15, -27, -19, 18, 10, -1, -16, -9, 29, 55, 31, 25, -24, 30, -24, -52, -19, -5, -41, -31, -12, -3, 10, -21, -2, -20, -9, 15, 44, -21, -48, -38, -10, -27, 37, -12, 0, -3, 0, 22, 41, -1, -39, -2, -24, 13, 26, -32, 36, -7, -15, 14, 24, 5, 7, -35, 10, -32, -26, -27, 14, 3, -30, -19, -28, -24, 20, 20, -36, -29, 2, -27, -3, -19, 31, 46, 23, 13, -14, 5, 8, 26, -1, 34, 19, -18, 28, -39, 10, 30, -44, 9, 26, -24, 36, -25, 3, 20, 36, 53, 37, 15, -25, 14, -16, -30, -22, 1, -43, -11, -35, 12, 32, -6, 23, -41, 13, -6, 25, 17, -15, 17, -30, 46, -12, 38, -6, 10, 10, 17, 0, -38, 4, -14, 21, 11, 34, -19, 4, 18, 12},
  '{24, -10, 42, 6, 18, 1, -27, -8, 40, -3, -24, 30, -5, -17, -31, -18, -10, 27, 28, -35, 36, 18, -21, 3, 1, -20, -11, 3, 38, -27, -41, -26, 24, -3, 40, 9, -13, 47, 48, 46, 46, 19, 2, 38, -14, -3, 43, 43, -34, -19, -7, -29, -31, 17, -25, 11, 9, 63, 16, 15, 9, -16, -8, 39, 0, 12, 6, 37, 10, -20, -13, 16, 7, -2, -24, -5, 1, -9, -35, 11, 12, 22, 9, 22, -6, 8, 16, 23, 0, 5, -9, -17, 4, 20, 19, -11, -9, 15, 15, 57, 18, -35, 10, -31, -26, 41, 44, 48, 39, 26, -23, 8, 21, -11, 33, 23, -4, -2, -19, -32, 38, -33, 12, -25, 17, -34, 5, -28, -13, -16, -16, -32, 15, 4, 50, 5, 41, -6, 34, -15, 8, 26, 12, -16, -18, 18, -32, 16, -43, -12, -5, -21, 16, -19, 41, 27, 12, 39, 16, 29, 25, -16, 43, 7, -17, -21, -35, -43, -24, -47, -22, -34, 36, -46, -51, 4, -23, 13, 20, -19, 25, 40, 33, 44, 19, 29, 19, 6, 7, -5, 38, -24, -3, 5, -13, 29, -14, 29, 15, -41},
  '{-12, -10, -13, 23, 5, 14, -6, 16, -9, 26, -13, 43, -40, -48, -5, -27, -16, 14, -37, -11, -40, 14, 55, -15, 17, 1, 5, 53, 7, 6, -12, 16, 6, 93, 33, 36, 12, 7, 55, -16, -40, -58, -40, -6, -1, -13, 5, 11, -14, 34, -12, -27, 10, -31, -25, 13, -6, -28, -7, 11, 0, 30, -1, 11, 67, 1, 4, -17, -27, 27, 24, 50, -28, 10, 9, 21, 7, -29, -23, -39, -7, 7, -20, -26, -47, -16, 3, 11, -7, -11, -20, 43, -9, -12, -13, -30, 1, 27, -7, -30, -19, 1, 15, -19, -38, -1, 27, 47, -34, -12, 42, 11, 9, 6, 33, 17, -8, 2, 3, -3, 23, 32, -27, 0, 0, 28, 12, 28, 1, 7, 8, 10, 43, 44, 8, 6, -11, -14, -7, 3, 19, -19, 17, 10, 19, 14, 31, -5, 3, -8, 7, -31, 3, -15, -15, -7, 17, 22, -12, -35, 10, 4, 5, -35, 32, -8, 31, 14, -21, -16, 21, 34, 45, 24, 41, 15, 21, 13, 32, -6, 4, -14, 12, 40, 21, 25, 37, 15, -44, -11, -30, 36, 1, -13, 41, 6, -4, -5, 10, -1},
  '{-39, 1, -54, -52, -21, -21, 7, -35, 17, 38, 22, 8, -24, 17, 7, -31, 20, 5, -15, 10, -50, -2, 4, 0, -27, -29, -66, -45, 12, 35, -23, -76, -62, 6, 38, -78, -38, -27, 17, -12, -30, 13, -11, -22, -32, -5, 40, 11, 45, 32, -15, -19, 31, 33, -23, 33, 41, 1, -12, -19, -17, 2, -70, 39, 33, 34, 45, -17, 48, 36, -6, 24, 10, 27, -8, 47, -12, 30, 17, 35, 17, 10, -12, -1, 27, -23, 32, -15, 32, -30, -31, -8, 0, 9, 7, -29, 31, 2, -22, -9, 8, 6, 1, 18, -39, -1, 15, -25, 11, -22, 27, 46, 13, -44, 0, -2, 22, 26, -12, 15, 29, -9, 14, 23, -34, 6, -7, -18, 13, 39, -45, -34, -71, -18, -10, -31, 10, 16, 9, 36, -18, -18, -44, -10, 48, -28, 27, 30, 32, 28, -1, 9, -1, -13, 14, 6, 19, 10, -42, 12, 34, -11, 18, -39, 38, 24, 32, -32, 39, -11, -12, -22, 20, 6, -16, -23, 38, -3, -35, 33, -13, -24, 22, -18, -19, 4, 42, -28, 6, -10, -6, 9, -31, 28, 10, -25, -17, 42, -9, 0},
  '{-6, 40, 1, 37, 37, 13, 13, 1, -27, 18, 18, 39, 23, 20, 15, 8, 39, -29, 32, 14, 59, 7, -35, -10, -12, 25, -1, 3, 61, 55, -10, 50, 55, -32, 0, -9, 21, 3, -15, 15, -4, 57, 52, 44, 44, 69, 9, 23, 5, 16, -20, 29, -11, 15, 12, -10, -13, 25, 24, -46, -27, -31, 21, 43, -5, 14, 3, 15, 17, 26, -8, 13, 23, 27, 11, -19, 22, -36, 40, 2, 1, 10, -25, 10, 3, 9, 11, 27, 30, -40, 28, -37, -8, -12, -38, -13, 19, 5, -13, 18, 17, 41, -27, -39, -26, -15, 0, -4, 4, 32, 24, 15, -26, 26, 46, -35, -22, 18, 52, 32, -35, -26, -14, 3, 9, 28, -10, -29, -13, 7, 40, 48, -2, -17, -29, -23, 50, 1, -11, -41, 56, 16, 14, -12, 11, -20, 20, -7, 42, 1, 17, 16, 22, -24, 15, 30, 29, -30, 8, -11, -13, 26, -8, -12, 27, 27, -14, 19, -5, -21, -37, 6, -7, -3, -8, 12, 30, -10, -5, 25, 32, 23, 40, 39, -26, 0, 0, -6, 51, 20, -28, -26, 39, 22, 36, -20, -11, -33, 13, -29},
  '{21, 45, -25, 26, 16, 11, 28, 14, 10, -24, 61, -37, -50, -11, 13, 0, 13, 29, -25, -1, -11, 8, -35, 45, 8, 20, 48, 18, -31, -22, 62, 89, 14, -59, -86, 49, 7, 38, 16, -60, 22, -23, -49, 40, 37, -51, -46, -19, -18, 46, 8, 27, 59, 35, -13, 11, -21, 5, 22, -26, -24, -34, -11, 9, -26, 29, -6, -4, -23, -13, -13, -23, 12, 18, 24, -26, -25, -14, 9, -26, -24, -24, 22, 14, 34, 20, -39, 7, 44, 40, 1, -4, 36, 18, -6, 13, 26, -8, -2, -32, 11, 12, 16, -12, -21, 7, -15, 3, 48, 40, -1, 1, 39, 11, -1, -23, 3, 42, 24, -32, 8, -4, -1, 18, 9, 16, 29, 29, -36, -39, -1, 49, 49, 5, -4, 9, -48, -8, -7, -13, -12, -42, -39, 24, -5, 14, -15, 30, -20, 2, -5, 1, -23, -4, -21, -10, -15, -12, 26, 24, 20, -27, 29, -15, -27, 28, 24, 48, -3, 17, 18, 4, -21, 25, 33, 27, 21, 3, 36, 28, 22, -28, -20, 38, 10, 39, -43, 27, 29, -24, -10, 23, -4, -6, 9, 33, -5, 36, 2, 27},
  '{0, 0, -1, -6, -3, 3, 1, 3, 13, 9, -2, -1, -3, -1, 11, -11, -8, -9, 1, 2, -2, -4, 8, -1, 1, 1, 1, 1, 0, 0, -1, -1, -1, -1, 0, 1, 1, -13, 13, 12, 0, 1, 1, 4, -1, 0, -7, 7, 2, 1, -1, 0, -3, 1, -1, 1, -10, -7, -2, 0, 1, -1, 3, 12, 7, 7, -3, 0, -3, 0, -2, -2, -2, 1, 1, 0, -1, -2, -1, -1, 1, -9, -1, -1, -1, 2, -2, 0, -2, 3, -4, 16, 0, 2, 2, -3, -15, 0, 3, 1, 0, -1, -3, 0, -3, 1, -1, 11, -3, -14, 1, -3, -2, -3, -6, -4, -8, -9, -4, 1, -1, 7, -9, -1, 1, -1, 1, 0, 0, 0, 1, 0, -1, -2, -1, 1, -7, -1, -8, 6, 0, -3, -6, 2, -8, -5, 11, -5, -1, 1, 0, 0, 0, -5, -2, 1, 5, 18, -1, 4, 1, -1, 8, 13, -1, 7, -1, -2, -9, 0, -1, -2, 13, 1, 2, 0, -2, -2, -3, -2, 1, -6, -13, -15, -5, 0, -9, -1, 3, 6, -11, 6, -6, -1, 0, -13, -4, -15, 0, 1},
  '{10, -2, 16, -12, -23, -11, -3, -12, -2, 20, 15, 6, 26, -10, 14, -8, -13, 21, -17, -4, -26, 26, -9, 0, 49, -9, -29, 10, 38, 7, -2, -16, 30, 14, 45, 23, 5, -2, -21, -65, -8, 26, -6, 10, 3, -12, -11, -3, 26, -5, 15, 16, -2, -5, 11, -15, 39, -21, -13, 11, 11, 5, -13, 22, 3, 14, -18, 1, 15, 8, -13, 9, -6, 30, 35, 21, 22, 35, 4, 9, 11, 15, 7, -16, -18, 6, 6, -11, 15, -7, 6, -27, -17, 32, -18, -5, -5, 12, 19, -8, 48, 26, 6, 35, 12, -2, 10, 24, -26, -10, -11, -20, -46, 12, -32, 11, -27, -17, 10, 11, 27, 18, -12, 22, 18, 22, -3, -20, 25, 16, 5, -9, 26, 42, -12, -17, -7, 4, 1, -31, 13, -10, -28, -5, 9, 8, -1, 2, 4, 29, 26, 28, -1, -4, -8, -6, 32, -11, -29, -34, 0, -38, -27, -4, -32, -9, -26, 6, 10, 11, 19, 0, 3, 32, 25, 42, -9, -1, 10, 27, 10, -19, -13, 18, 4, -26, 3, 12, -41, 36, -17, -34, -2, 0, 39, 15, 13, 8, -26, 39},
  '{22, -7, -24, -34, -12, 28, 33, 11, 41, 2, 9, -27, 29, 26, 36, 1, -12, 12, 45, -1, -65, -52, -45, 31, -35, 4, -17, -5, 36, 48, -9, -58, -59, -31, 51, 29, -25, 20, 17, -12, 54, -36, -11, 15, 45, -8, -29, -15, -8, -26, -17, -5, -3, 34, 37, -17, 23, -23, -34, -6, 47, 0, 47, -3, -9, 27, 30, 16, -16, 20, -14, -6, 41, -22, -34, 40, 18, 25, 16, 71, -16, -6, 42, 37, 29, 47, 3, -8, 0, 0, 32, 9, 41, 5, 23, -10, 48, 30, -11, 4, -6, 0, -1, -22, -6, 19, 33, -22, -4, 31, 23, -26, 25, 29, -4, -27, 25, 23, 33, 7, 19, 3, -28, 26, 21, 8, -47, -2, -18, 9, 9, -24, -60, -3, -13, 19, -23, -20, 6, 25, -16, 20, -4, -5, 37, 2, -6, 8, -19, -33, -19, 16, 14, -33, 30, -22, 33, 20, 11, -23, -9, 8, 32, 3, 16, -34, 4, 49, 45, 31, -37, -40, -18, -34, 7, 14, 12, -30, -36, -9, -11, 11, -19, -11, 7, -10, 15, 22, -1, -21, -24, 15, 33, 1, -25, -4, -32, 39, -15, -1},
  '{23, -6, 15, 41, -31, 13, -33, 42, 14, -25, 5, -13, 1, 13, 28, 28, 10, 9, 36, -2, 0, -27, 46, 17, -2, -17, -37, -28, 49, 74, 17, -48, -36, 26, 3, 52, 21, -36, 15, 41, 29, -29, 24, 10, -9, -29, 31, 5, -54, -28, 34, 29, -8, 5, 26, 41, -21, 4, -48, -5, 35, 52, 42, -7, 25, 10, -26, 19, -4, 5, 19, -2, -24, 4, 11, -14, 12, 32, -1, 6, 12, 34, 18, -44, 1, 30, 11, -20, -48, -32, 8, 28, 44, -22, 17, 8, 38, -14, -8, 1, -31, -23, 40, -26, -22, 9, 0, 42, 9, -41, 8, 31, -7, 10, 2, 18, 22, 33, 19, -47, 34, 20, -7, 18, -10, 23, -29, 16, 35, 34, -22, -4, -28, 5, 31, -11, 9, 22, -3, 51, -16, -14, 41, 9, -39, -9, 19, -5, 10, -13, 32, 13, 39, 1, -31, 35, -2, -5, -8, 17, 8, -8, 24, -3, -38, -11, -17, 28, -19, 22, -16, -28, 18, 9, 27, -25, 37, 31, 30, -17, 1, 16, -5, -35, -27, -28, -8, -2, 3, -43, 9, -15, 0, 34, 18, 35, 35, -16, 46, -7},
  '{37, 33, 20, -34, 33, 38, 12, 0, 41, 35, -26, -41, -7, 29, 3, 39, 28, -29, -3, 40, 9, 23, 17, -13, -14, -23, -12, 57, 20, 12, -2, 59, 22, 17, 40, 10, 4, -17, 48, 42, 26, 71, -2, 1, -26, 57, -7, 9, 33, 38, 14, -29, -42, -11, 9, 37, -6, -24, -46, 24, -32, -37, -4, 16, 28, -5, -22, 32, 38, -11, -11, 1, -7, -4, 5, -8, 16, -44, -1, -2, -30, 7, 0, -39, -8, -18, 26, 43, 0, -59, 8, 5, 14, -11, -7, 12, -2, -20, 1, -9, 48, -24, -7, 10, -34, -6, 0, 15, 19, 19, -28, -18, 12, -33, 29, -17, -6, -20, -10, 42, 19, -30, -2, 19, -6, 20, 45, 6, -12, 34, 27, 19, 21, 15, 53, 28, -31, -24, 19, 30, 4, 3, -19, -21, -27, 4, 4, -7, -12, 13, 20, 41, -36, -36, 12, 7, 8, 1, 38, 13, -28, 24, -2, 23, -13, 0, -37, -47, -27, 18, -9, 26, 11, -6, 0, -15, 35, -18, -28, -7, -1, -12, -5, 42, -16, -9, -20, 25, -1, 19, 29, -25, 4, -5, 19, -26, 35, 41, 15, 15},
  '{27, 14, 8, 14, 37, -13, 32, -7, 29, -13, 1, -1, -2, -25, -42, 50, 21, 7, -3, 26, 3, 50, 46, 36, 12, 30, 42, 39, -61, -61, 48, 33, 33, -50, -64, 29, 13, -40, 1, 91, 30, 11, 5, -12, 23, 19, 16, -58, -43, -24, -31, 15, 10, 13, 9, -20, 37, 29, -4, -27, 8, 52, 6, -2, -4, -14, 5, 40, -14, 37, -12, -44, -2, 4, -3, -8, -4, -14, 11, -56, -9, 7, 0, 16, 7, -10, 8, -4, -21, -40, 7, -8, 15, -46, 6, -1, 15, -14, -28, 7, 14, -9, 59, 55, 5, -35, -47, 7, -27, 35, 20, 24, -3, 38, 4, -27, -10, 30, 9, -30, 56, 23, 40, -3, 52, -2, 13, 39, 21, -46, 51, 46, -6, -14, -30, -24, 17, -2, 41, 32, -44, -14, 35, 27, -40, 1, 11, 10, 29, 46, -21, 3, 2, -15, 26, -2, -50, -19, -19, -13, -13, 4, 46, 12, 10, -7, -6, -27, 8, 29, 18, 34, 14, 39, 63, 7, 13, 19, 4, 50, 0, 4, -18, 1, 4, 6, -16, 50, -2, 12, 10, -35, -1, -11, -33, 13, 0, -14, 25, 32},
  '{-13, -27, -11, 13, 28, 30, 13, -16, 17, 28, -2, 11, 39, 46, 13, -16, 38, 5, -7, -33, -1, -53, -16, -27, -30, -38, -55, 7, 4, 37, -5, -68, -58, 0, 6, -73, -73, -33, -70, -12, 20, -28, -23, -25, 12, 24, -38, 25, -38, -9, 29, 34, 31, 29, 14, 8, 46, -1, 17, 14, -3, -30, 22, 5, -32, 39, 43, 26, -11, 10, -20, 28, 55, -4, -29, 13, 29, 51, 54, 45, 33, 26, 36, 44, 20, 24, 3, -12, -7, 41, 9, -4, -6, -4, -6, 21, -2, -3, -3, -15, 39, 37, 13, 6, -27, 2, 20, -32, -16, -11, 23, 28, -3, 53, 45, 13, 8, -16, 38, 3, 1, 24, -31, 14, -37, 24, -8, -3, 3, 36, -5, -7, -32, -64, -24, -32, -12, -39, 10, 24, 22, -3, -1, -13, 24, -48, 2, -25, 1, -31, -27, 37, 41, 29, -33, -15, 44, 31, -35, 15, 30, 19, 14, -19, 27, 2, 6, -26, -14, 19, -32, 4, -17, -22, 1, 41, 33, -30, 19, 7, -20, 14, 35, -23, 35, 23, 11, -4, 11, 30, -10, -15, -22, 19, 13, 13, -43, -10, 3, -26},
  '{17, 0, -15, 2, 26, -16, -12, -29, 18, -47, 27, 6, 30, 0, -6, 23, 12, 19, 10, 19, 18, -5, 55, 29, 11, 29, 21, -29, 6, 62, 40, 6, 23, -1, 21, 44, -21, -55, 53, 37, 16, -35, -39, 7, -11, -35, 11, 22, 19, 7, 3, 32, 2, 41, 3, 35, -9, -30, -19, -21, 15, -13, -41, -36, 60, 4, 24, -38, -47, 27, -20, 12, 22, 36, 19, -1, 32, 30, 58, 68, -9, 16, 44, 4, 41, 29, 0, 29, -10, -6, -25, 0, 28, -13, -25, -23, -4, -31, -45, 0, -21, 33, 11, 48, -19, 10, -37, 4, -18, 18, 4, 27, 43, 26, 8, -20, 40, 49, 36, 22, 2, -8, 56, 47, 59, 17, 5, -17, 45, 41, 44, 4, -1, -6, -8, -4, -8, -24, -25, 31, 15, 15, -21, -19, -5, 3, 37, 58, -2, 9, 31, 13, 16, -4, -34, 16, -20, 32, -53, -35, 37, 25, 33, -47, -26, 16, 9, 24, -29, 9, 36, 12, 48, 18, 33, -19, -24, 20, 10, -29, 8, -34, -19, -15, -27, -35, 21, -1, -13, 33, 18, 58, -14, -36, 9, -17, 14, 13, 0, 43},
  '{-31, -26, -1, 21, 12, 29, -19, -8, -8, 20, -13, -9, 36, 6, 52, -16, 6, 17, -33, -12, 1, 20, 24, -38, -58, 21, 17, -31, -47, -75, -37, -18, -53, -60, -44, -51, -69, -5, -22, -9, -11, 14, -34, 8, -11, 35, 17, -2, -14, -47, -9, 1, 17, 19, -2, -3, 11, -23, 10, -23, 2, -27, -54, 18, -16, 18, -7, -1, 4, 16, 0, 10, 20, 5, -1, 20, -17, 38, 4, 2, -14, 43, 11, 26, 21, 11, 7, -18, 27, 32, -17, 1, -24, 26, 33, -45, 12, 9, -4, 4, 12, -3, 10, -26, -2, 4, 1, -2, -13, 10, 1, 39, 22, -11, -3, 26, -6, -44, -15, 17, 15, 18, -36, 39, 14, -8, -16, -8, -35, -24, -26, -48, -44, 34, -31, -47, -6, 0, -9, -22, 39, 47, 33, -2, 13, 10, 29, -24, 4, -28, 3, 15, 36, 10, -11, -12, -14, -14, -25, -11, -17, 11, -10, 35, 44, -15, -38, -26, -18, 45, 24, -29, 10, 39, 14, 1, -29, -1, 9, -16, 18, 38, 24, 38, 54, 43, 34, 10, 32, 43, -4, 9, 12, 35, 47, 5, -19, -18, 29, -19},
  '{10, 33, 25, 34, -16, 14, 14, -17, 51, 30, -26, -35, -7, -3, 26, -3, 1, -35, -11, -40, -4, -40, -37, -45, 0, -19, 66, -16, 12, 9, -27, -10, 69, 25, -54, 21, 15, 46, -31, 2, 4, 4, -11, 0, 13, -27, -4, -14, 7, -45, 22, -47, -42, -47, 0, 2, -29, 7, 62, -7, 27, -22, -8, -1, -1, 40, -15, -27, 17, -34, -37, 10, 42, -2, 34, -42, -20, -21, -37, -26, -12, -4, -45, -14, -20, 37, -16, -7, 6, 43, 33, -5, 17, 14, -8, 18, -30, -9, 11, 7, -25, 24, 23, 24, -38, 4, -10, 21, -13, -4, 12, -40, -39, 18, 29, -38, -22, -3, 50, 25, -22, -32, 21, -22, -4, -36, -3, -30, -12, -15, 17, 14, 54, 43, -15, 16, 15, 23, 32, -21, -23, -2, -8, 29, -44, 5, -42, -23, -42, -45, -32, -16, -9, -20, 34, 2, -12, 11, -13, 35, -35, -43, -18, 40, 7, -20, 17, 52, 25, -31, -13, 13, -16, 3, -40, -38, -41, -11, -4, 25, 9, 21, 0, 49, 39, 8, 17, -1, 6, -23, 22, -41, -22, 35, 12, 2, 9, -9, 31, -45},
  '{2, -21, 5, -2, 14, -9, 38, -21, 35, -13, 14, 0, 33, 36, 12, 58, -3, -24, 29, -13, 15, 38, 60, 30, -6, 16, 30, -9, -12, -70, -17, 35, 26, 11, -70, -6, 1, -17, 19, 28, 24, 0, 34, -5, -46, -7, -6, -1, 18, -6, 13, -42, -34, 0, 5, -39, -35, 52, 41, 7, 11, -29, -18, -54, 24, -20, 17, 14, 1, 27, -12, -2, 21, -34, -17, 0, -11, 25, -9, -54, 26, -23, -39, -24, -10, -28, -15, 9, -45, 23, -36, -3, -29, -18, 8, -37, -40, -46, -8, -3, 32, 30, 44, 9, -13, -12, -37, -16, 14, 45, -44, -6, 34, 24, 7, -13, 11, -16, 8, 39, 5, -20, -28, 44, -12, -35, -5, 62, 19, -30, -8, 28, 34, 20, 21, 17, 8, 8, 19, 34, -28, 28, 4, 18, 1, -5, -26, -33, 16, -9, -1, 4, -9, -1, 9, 29, -2, -31, -8, 9, -6, -12, 8, -16, 18, 5, -18, -1, 18, -2, 45, -5, -14, 39, 40, 7, -12, 49, -5, 29, 29, -32, 31, 12, 40, -9, -12, 14, 15, -10, 36, -15, -40, -14, -25, 35, 27, -10, 2, 34},
  '{-29, 3, -23, 23, 32, -43, 12, 12, 14, -27, -11, -5, 38, 26, 34, 5, 23, 19, 15, 35, -68, -23, -20, -18, -5, 17, -4, -15, 51, -6, -49, -109, -56, 1, 56, -3, -67, -9, 2, -4, -31, 11, 12, -5, -9, 33, -14, -32, -23, 27, 9, 1, -25, -7, -28, 22, 25, -31, -36, 34, -22, -2, 13, 2, 54, 45, -9, 9, -8, 41, 16, 36, 27, 25, 12, 17, -5, 13, 18, 71, -4, 12, -8, 33, 48, 17, 42, -23, 19, 3, -11, 37, 6, 9, -23, 11, 3, 2, 12, -23, 28, -16, 30, -2, 33, -26, 17, -35, -47, 22, 14, 38, -22, -2, -24, 9, 24, -17, 34, 27, -26, 35, 5, -28, -26, -27, -53, -39, -20, 32, -35, -2, -23, -17, 10, -15, 4, -21, 2, 0, 30, -27, 17, 11, 42, -23, 2, 14, 8, -6, 8, 22, 33, 2, 18, -13, 46, 0, -1, -31, 3, 0, -24, -34, 28, 36, 43, 15, 42, -25, 19, 15, 4, 41, -11, -23, -17, -37, -9, 6, 18, -10, 26, 9, -26, 38, 48, -9, -42, 17, 6, 43, -5, -22, -24, -22, -19, 30, 2, -27},
  '{-13, -13, -17, 5, -38, 23, 40, 24, -3, 33, -1, 13, 3, 26, -28, 23, 27, -13, -25, -15, 1, -20, 7, 12, -9, -6, -9, 8, 21, 31, 4, 8, 25, 22, 12, -6, -18, -22, 2, 24, 10, 3, 27, -28, -25, 22, -7, -5, -23, 3, 10, 2, -41, -33, -24, 25, 8, 5, -3, -6, 19, 10, 15, -18, 29, -15, 2, 0, 11, -1, -21, 8, 15, 0, 11, 7, 6, -26, -35, -21, 4, 8, -33, -28, -11, 3, 16, -3, -14, -13, 9, 14, -17, 6, 23, -7, -1, 2, 20, 19, 1, 14, 14, -32, 13, -17, 24, -7, 11, -4, 10, 28, 1, 0, -4, -5, 36, -7, -19, -28, 1, -5, -2, -6, 37, -1, 1, 5, 13, 11, 12, 14, 0, 2, 7, -8, 0, -9, 10, 9, 14, 13, 0, 2, -1, -4, 3, -9, -6, -2, -22, 22, -10, -19, -33, -20, -2, -6, 4, 0, -4, 13, -25, -12, -29, 16, 38, -27, -33, 27, 3, -14, -1, -12, -4, 21, -10, 3, 5, -14, 31, 9, -9, -15, 25, -2, 12, -1, 6, 19, -29, 0, 18, 8, 30, -14, -17, 17, -22, 38},
  '{-21, 26, -23, -11, 33, 24, -7, 31, 56, -29, -15, -34, -29, 5, -56, 38, -31, 6, 27, -20, -35, -3, 26, -25, 46, 50, 50, 24, 9, -64, 1, 7, 67, 14, -73, 29, 59, 37, -1, -25, -5, 10, -11, 18, 17, 19, -53, 5, -2, 5, -5, 1, -1, 5, -2, -22, 4, 16, 23, 23, -4, 24, -7, 4, 4, 10, 18, -46, -60, -14, -34, -10, -27, 31, 43, 4, -6, -33, 14, -21, -19, -37, -7, 22, -2, -2, -38, 21, 3, 27, -8, 16, 22, 11, 1, -18, 8, -26, 4, -2, -31, -4, -1, 28, -28, 14, 9, 35, 39, 45, 15, -48, -19, 44, 34, -24, 14, 1, 40, -41, 20, -24, 3, 15, -22, 32, 14, 35, 16, -33, -9, 45, 29, 54, -13, 48, 30, -21, 16, 21, -37, 4, -42, 27, 7, -41, -19, -11, -25, -10, 5, 30, 32, 4, -9, 28, -19, -17, 31, -22, -15, -7, 10, 12, 10, -19, -11, 32, 12, -13, 23, 28, 11, -21, -16, -1, -23, 16, -4, -13, -33, -9, 4, -10, 45, 6, -9, 0, -23, 1, 8, 7, 40, 25, -4, 3, -32, 29, -9, 10},
  '{15, 28, 6, 10, 49, 34, 6, -8, -4, 5, -5, 11, -21, -34, 29, 5, -38, -30, -12, 1, -15, -12, 30, 4, -36, 14, 26, -31, -20, -82, 9, 3, -3, -37, -84, 1, -45, -37, -19, 19, 17, 7, -20, 5, -4, -36, -16, -24, -34, -28, -37, -35, 22, 10, -2, 34, 43, -14, 28, -42, 19, 6, 24, 24, 12, 37, -20, 17, 26, 20, -3, -3, 6, -25, 5, -4, -14, 0, -9, 12, 14, 9, 29, -1, 29, -22, -25, -20, 11, 3, 4, 28, -7, 11, -31, 2, 11, 21, 4, 24, 25, -18, -15, -28, 46, -8, 21, 2, 30, 10, 40, 43, 42, 0, 22, 45, 1, -4, -18, -25, -28, 29, 16, 35, 4, -44, -35, -4, -17, -21, 7, 7, -32, 17, -18, -6, 34, -25, 13, 31, 16, 33, -7, 28, -2, 20, -27, -35, -9, -17, 12, 40, 10, 39, 2, 24, 39, 12, -24, 34, -23, 26, -20, -13, -15, 14, -18, -22, 1, 15, -17, -24, -20, -7, 1, -10, 40, 25, -27, -2, 27, -33, -16, 27, -11, -22, -29, -4, -8, 29, 10, 21, -16, 31, 13, -22, -32, -35, 28, -30},
  '{33, -30, -20, 30, -25, -34, 29, -20, 22, 4, 29, 23, 28, 34, 42, 35, 46, 46, -18, -21, -12, -5, -11, -3, 15, -7, 42, -23, 4, 44, -30, -9, 54, 13, 33, -45, 19, -32, 8, -25, -4, 18, 33, -39, -29, 29, 68, 50, 33, -4, -36, -9, -23, -16, -18, -33, -17, 9, 25, 23, 12, 24, -5, 51, 5, 6, -23, 37, 8, 7, 14, 7, 20, -15, 23, -10, -36, -20, -40, -12, 11, 35, 4, -22, -49, 0, 32, -3, -19, 0, -37, -14, -25, 13, 0, -37, -10, -26, 11, -17, -36, 16, -13, 11, -4, -31, 33, -33, 9, -19, -6, 34, -39, -22, 12, -24, 23, -20, 6, 46, 5, 14, -3, -14, -2, -24, -22, 26, 33, 7, 10, 2, -33, 37, -16, -13, 10, 9, 28, -3, 25, 46, 26, -5, 16, 27, 22, -7, 27, 2, -37, 20, -4, 30, -5, 25, 31, -14, 7, -19, -24, 25, 27, 18, 10, 6, -14, -31, -7, -21, 16, 43, 19, 0, 28, 25, 26, 46, 1, 16, 0, -25, -31, -10, 38, 29, -12, 18, -13, 25, -16, 1, 7, -9, 28, 15, -26, -3, -18, -9},
  '{0, -20, -32, -6, 27, -19, -8, -21, 2, -17, 2, 29, 21, 28, 0, 42, 29, 42, 30, -1, -22, 25, 31, 40, 63, 37, 13, -15, 41, 73, -63, -14, -34, 70, 87, 49, -12, -6, 11, 71, 29, -67, 1, 1, -75, -25, 29, -33, -43, -29, 14, -11, -13, -21, -39, 43, 11, 39, -48, 23, 37, 38, 19, -52, 80, 29, 8, 19, 38, -4, 41, 26, -5, 37, -16, 5, 16, 16, 18, -13, 39, 24, -13, -26, -51, 25, -8, 24, -55, -30, 0, -19, 8, -26, 3, 32, 31, -24, 3, 27, -25, 13, 54, 23, 19, 13, -26, 36, 10, 6, 6, 26, 27, 23, -21, -18, 17, -9, -32, 17, -17, 16, 7, 54, 35, 13, 9, 18, 26, 80, 11, -19, -22, 18, 32, -15, 20, 19, 3, 34, 3, -31, -3, 15, -35, 28, 49, 19, 32, 1, 13, 13, 57, -6, -16, 14, -38, -18, -24, 3, -42, 10, 30, -25, -8, -16, 22, -21, 22, -20, 38, 42, 43, 27, 66, -39, 43, 0, -7, 43, -1, -37, -13, -8, -1, -35, 3, 21, -3, -36, -42, -12, 22, -2, 21, 32, 41, 11, -4, -5},
  '{-44, -15, 47, 27, 15, 2, -15, 9, 18, 37, 26, 6, 42, -19, -25, 4, -18, 15, -6, 0, -4, 6, -14, -17, 60, 20, 31, -35, -34, -1, 25, -49, 15, -11, -18, 19, 31, -50, -15, -28, -8, -80, -19, 22, 25, 0, -13, -42, -22, -3, -11, -19, 34, 24, 15, -28, -11, 12, 15, 38, 39, -10, 24, -12, 11, 14, -30, -21, 2, 15, 11, 13, -35, 31, 21, 22, 0, 33, -28, -43, -29, 29, -27, 1, 2, 33, -30, -9, 17, 63, 4, -9, 10, 0, 29, 11, 5, -7, -5, 20, -34, 16, -17, -11, 45, 27, 26, 10, 25, 38, 11, 33, 7, -21, 32, -6, 37, 38, 11, -10, 38, 44, 23, 2, 43, -18, -9, 42, 7, 1, 14, 11, 0, 27, -43, 26, -26, -37, -14, 13, -46, -2, -14, 10, -6, 7, 2, -36, -42, 33, 13, -2, 11, 0, -22, 12, -29, -15, -37, 22, 21, 29, -18, -29, -16, -11, 47, 34, 24, -16, -8, 25, 18, -19, 25, -2, -34, -19, -15, -10, -12, 24, -29, 7, -9, 15, -22, -22, -32, -1, -21, 42, 10, -14, 12, 35, 20, 18, -15, -14},
  '{-38, -4, -23, 15, 13, 6, 33, -21, -30, -27, -10, -15, -18, 33, -12, -12, 4, -9, -32, -15, -3, 41, 42, -18, 36, -6, -35, 13, 74, 69, -49, -36, 17, 22, 69, -48, -53, 17, 4, 22, 23, 32, -11, 13, -42, 19, 7, 57, 50, 0, 6, 23, 26, -40, -10, -28, 8, 6, -13, -6, -26, 28, -22, -7, 34, -18, 25, -26, -6, 3, -26, -5, -4, -9, 18, 7, -12, 4, 33, 18, 10, 20, 15, -11, 5, -16, 18, -3, -2, -51, -23, 2, -3, 41, 41, -33, -8, 5, 15, -3, -8, 5, 1, -24, 0, -36, -2, 10, -33, 27, 36, 7, 16, -36, 0, 28, 1, 7, -21, -28, 8, 13, 33, 41, 2, 30, 11, -26, 29, 0, -49, -6, -2, 0, 40, -7, -2, 1, 12, 1, 8, 11, -18, 12, 2, 29, 10, 18, -14, 5, -7, 4, 21, -25, 23, 7, -2, 46, 12, -24, 28, -19, -33, -37, 2, -1, -16, -44, -22, -17, 2, -6, 30, 18, 45, 17, 23, 21, -8, 25, 11, -4, 22, -5, -23, -1, 44, 8, -26, 9, -2, 30, -10, -29, -10, -15, -9, -8, 29, -1},
  '{-24, -36, -33, 24, -11, 16, 6, -8, 17, 9, 49, 32, -13, 12, 18, 15, -26, 11, -11, 8, 15, -24, -33, -41, -34, 41, 27, 9, -5, -16, 49, -15, 23, 1, -56, -12, 12, 21, -40, -30, -6, 56, 23, 18, 62, -22, 28, 1, 49, 29, -12, -4, -12, 29, -9, -12, -5, 32, 3, -2, -21, 1, 4, 4, -50, -20, 6, 37, 20, 26, -15, -6, -9, -1, 43, 4, -35, -6, -25, 27, -16, -18, -8, 7, 11, 21, -4, -21, 21, 26, 38, 10, 1, 18, 7, 3, -16, 20, 4, -56, -4, 5, -32, -15, -11, -4, -28, 16, -11, -16, -17, 23, -19, -6, -10, -3, 4, 31, 3, -6, 7, -7, -21, -11, 8, -13, 1, 3, -5, -28, 9, 3, -8, -12, 6, -43, -1, 0, 11, -40, 16, 21, -12, 7, 17, -3, -8, 7, 10, -12, -8, -21, 13, -23, 8, -16, -2, 22, 19, -22, 32, 28, 40, -14, 17, -10, 21, -22, 28, 26, -2, -29, 13, 10, -36, 6, -2, 9, -22, -14, -8, -25, -19, -26, -41, 18, 47, 41, 35, -26, -8, 13, 22, -16, 20, -33, 16, -19, 2, -37},
  '{-49, 12, 15, 48, -8, 18, 40, -34, -27, 26, -29, 3, -17, -21, -13, -72, -13, -33, -19, -3, -9, -56, -14, -8, 2, -29, -26, -62, -61, 36, -16, -15, -46, -12, -22, -83, -85, -51, -28, -20, -44, -55, 7, -53, -34, -34, 10, -4, 14, -19, 25, 14, -14, 7, -18, 12, 21, 9, 44, 4, -14, -31, -34, 35, 10, 53, 16, -43, -19, -25, 27, 46, 27, -38, -22, -7, -4, -7, 12, -55, -18, 2, 3, -42, -20, -7, 24, 26, -1, 106, 2, 37, 7, 33, 40, -25, 59, -7, -19, -16, -38, -1, -3, 52, 12, 13, 47, -11, 42, 6, 32, 21, -19, 32, 44, 2, 17, 37, -11, 30, -44, 38, -12, 16, -29, 0, -11, 6, -9, 6, -35, -35, 31, -11, -23, -3, -25, 7, -12, -3, -20, 22, -6, 3, 11, -26, 1, 4, -12, 5, -10, -32, 4, 40, -3, 6, 13, 33, -17, 38, 45, -8, -7, -14, 43, 26, 30, -13, -21, -18, -15, 10, 1, -31, -11, -56, -40, 29, 43, -34, 31, 1, 5, 19, 11, 45, -19, 31, -29, 36, -20, -12, -29, 11, 17, 8, 30, -31, -22, -18},
  '{-9, -25, -11, -22, 4, 30, 30, 5, 26, 16, -8, 30, -11, -14, -31, -8, -5, 15, -30, -9, -5, -19, -29, -19, 9, -15, 19, 2, 5, -22, 1, -1, 0, 5, 4, -1, 8, 2, -26, 17, 9, 9, -9, 1, -1, 24, 13, -13, 0, 0, 1, 6, 5, 15, 8, -21, 1, 8, -11, -1, -12, -2, -28, 6, -10, 29, -6, 5, 9, -22, -22, 24, -26, -21, -3, 0, -9, -1, 15, -5, 0, -3, -3, 2, 0, 2, 0, -1, 1, 4, 1, 0, 1, 15, -6, -16, 2, 8, -13, -1, 6, 20, -14, 19, -13, -1, 12, 21, -38, 18, 5, -5, 13, -11, -5, -16, -34, -7, 0, 6, -4, -19, -1, -30, 26, 8, 6, -2, -1, -10, 0, -8, 14, -16, 9, 9, 26, 11, 3, -21, 10, -1, -3, 7, -8, 9, 9, -18, 2, -9, 4, -14, 3, 2, -2, -17, -38, -4, -25, 0, 18, 24, -21, -9, -11, 13, 15, 10, 1, -23, 17, 0, 10, -9, 21, -16, -17, -6, -23, 1, 31, -12, 33, -23, -2, 14, -21, 7, -16, -29, -2, -6, -21, -14, 1, -22, 23, -25, 14, 0},
  '{1, -36, 0, 28, 13, -1, -7, 1, -29, -5, 16, -16, -41, -64, -33, -17, 0, -9, -19, -5, 61, 39, 13, 16, 33, 12, 65, 39, -24, -20, 21, 39, 3, -57, -34, 46, 24, 16, 19, -5, -11, 15, 37, -10, 12, -4, -19, 28, 46, 17, -1, -29, 61, 6, 6, -25, 3, 39, 19, -8, -9, -7, -1, 2, -27, 10, -21, -16, -59, -8, 27, -37, 32, 28, 18, 22, -9, -17, -9, 7, -7, -9, 28, 20, 18, -14, -25, 0, 17, 31, -1, -16, -20, 2, 23, -17, -8, 5, 17, 6, 11, 3, -27, 50, 3, -24, -28, 28, 39, -2, 39, -29, -8, -3, -46, -3, -16, 21, 14, 30, 44, 19, 33, -3, 33, 13, 57, 10, -41, -9, 47, 34, 25, -23, -44, 22, -3, -20, 10, -8, -22, -28, -31, -34, -23, 17, 34, -16, 54, 42, -9, -10, -13, 0, -10, 9, 19, -9, -28, 24, -17, 9, 23, -46, -17, 19, -29, 33, -1, 3, 23, -22, 15, 26, 19, -24, 33, -30, 5, -10, -27, 13, 11, 41, -19, 21, -31, 11, -37, -15, 28, 39, 23, -4, 7, -13, 3, -11, 29, 50},
  '{44, -32, -22, -34, 22, -13, -33, -44, 1, -38, 17, 24, 35, 14, -35, -31, 3, 21, 20, 44, -53, -51, -28, 46, 6, -3, -8, -17, -51, -28, 40, -17, -40, -86, -21, 16, 20, -17, -41, 28, 10, -8, 5, -19, -3, -37, -26, -10, -17, 46, 20, 13, 14, 41, 45, 8, 26, -22, -32, -16, 18, 5, 2, -9, -29, 29, 17, 9, 10, -9, 12, 21, -18, 16, -10, -7, -8, 27, 67, 22, -27, -22, 18, 50, 85, -2, 21, -16, -2, 29, 5, 40, 56, -5, -27, 31, 37, -31, 4, -41, 22, 19, 39, -10, 30, -29, -20, 0, 16, -32, -3, -27, 40, 22, 10, -29, 21, 8, 2, 15, 12, 21, -13, -24, 23, -24, 28, 47, -1, 20, 32, 22, -21, -60, -46, -3, 24, 11, 15, -13, -8, -10, 34, 41, -7, -5, 37, 4, 29, -21, -13, 33, 35, -13, 27, -13, 20, -20, 18, 41, 28, 1, 43, 34, -1, 32, 1, 43, -4, -18, 24, -27, -30, -30, 14, 30, 13, -24, -5, 7, 31, -18, 30, 33, -31, -23, 16, 17, -19, -6, 28, 35, 46, 13, 17, 22, -26, 26, 18, -19},
  '{-34, 11, 18, -17, -22, -16, -20, 4, 3, -14, 21, 6, -58, -55, 12, 3, 24, -3, 3, -25, -3, -8, -2, -26, 11, -23, 9, -10, -15, -8, 15, 8, -6, 21, 2, -21, -30, 13, 36, -63, -42, 1, -12, 24, -17, -11, 21, 29, -6, 44, 30, 11, -20, 3, 16, 31, -1, 5, -22, 25, 11, 16, -27, 37, 44, 38, -1, 1, -26, 24, -2, 33, -4, -30, -24, 11, -15, 10, 15, 12, -20, 36, 34, 46, -10, -5, -27, 27, 33, 19, -26, 49, 16, 14, 32, 19, 32, -5, 3, -41, -27, 30, 6, 36, -20, 35, -9, 24, 30, -8, 19, -1, -17, 9, 7, -22, 37, 23, 32, 5, -16, 48, 35, -5, 47, 0, -11, 18, -6, 29, -1, -4, 28, 42, -14, -29, -50, -26, 1, -7, 23, -44, -39, -41, 43, 5, -22, 3, 30, 14, -3, -36, 6, 17, -28, 2, 1, 33, -31, -2, 4, 21, -44, -25, 9, 10, 23, 19, 40, 20, -28, 37, 47, -30, -24, -26, -15, -31, -25, -39, -4, 28, -29, 36, 6, 27, 21, -43, -40, 43, 37, 55, 29, -5, 28, -40, -24, 45, -28, -11},
  '{-26, -39, 30, -8, 23, -25, -5, 2, 40, 31, -2, 23, 53, 39, 26, -10, -6, -15, 12, -44, 2, 35, 11, 24, -38, -19, 28, -58, 7, 9, -15, -99, -40, -27, 64, -35, -10, -18, 32, 35, -11, -2, 44, 0, -15, 12, 22, -21, -17, -10, -31, 25, -19, -27, -64, 7, -32, 18, 22, 40, 29, 51, 23, 4, 51, -35, -9, 15, 7, 4, -5, -14, -2, -1, -53, -45, -20, 30, 21, -8, -11, -21, 21, -54, -23, -28, 30, -11, -63, -22, -31, -8, -15, -31, -16, 19, 15, 20, -2, 16, -20, 2, 35, -2, 31, -42, -21, 42, -30, -30, 8, -29, -6, 5, -38, 16, -24, 2, 17, -13, -2, 22, 33, 39, 29, -25, -36, -59, -20, 58, -45, -15, 7, -1, 4, 3, 18, 38, -1, 49, -29, 3, 1, 18, -55, -23, 26, -16, -33, -30, 4, 16, -15, -3, 36, 25, -21, 0, -11, -31, -41, 20, 12, 46, -3, -9, -38, -26, 9, -9, -40, -8, 41, -20, 2, -22, -39, 8, 20, -27, -36, 4, -7, 15, -3, -12, -30, 38, -19, 6, -1, 25, -4, 0, -54, -32, 21, 35, 19, -30},
  '{-24, 9, 0, -12, 19, 20, -34, -23, 20, 37, 6, -14, 19, -6, 45, 37, -3, 39, 12, 33, -40, -15, 26, -14, -14, 26, -8, 11, 11, 26, -20, -29, 13, 17, 19, -64, -54, -8, 45, 24, 15, -29, -41, 21, 45, -13, -22, 7, -26, -14, -12, 18, 22, -5, 17, -25, -1, -36, 8, -25, 18, -5, 14, -1, 7, 34, 1, 12, 22, 13, -18, 22, 36, -31, -20, 5, 6, 33, 12, 37, -27, -12, 13, -13, 10, -6, 30, -5, -29, -23, -7, -23, -18, 41, -32, -7, -22, 41, 10, 27, 31, -9, -4, 10, -18, -4, 4, 2, -11, 8, 23, 22, -40, 9, 38, 15, 8, -19, -10, 7, 10, -8, -32, 23, 12, 19, -59, -2, -22, -3, -21, -30, 14, 2, 59, -32, 34, -9, -15, -6, 10, 9, -11, -4, 35, 7, 9, 12, 5, 12, -20, -1, 21, 13, 42, -11, 4, 34, 24, -2, -23, -3, -29, -2, 8, 14, 22, -34, 2, 40, -21, -24, -4, 32, 12, -24, 32, -47, 14, 23, 8, 52, -17, -24, 12, 29, -7, 7, 10, -8, -9, 18, -6, 19, 0, 3, 23, 5, 10, -21},
  '{40, -3, -26, -18, 5, -10, -21, 22, 3, 18, 37, 6, -13, 32, 17, 44, -2, 15, 39, -4, 25, -48, -31, -19, 68, 51, 25, 18, 47, -6, 84, 28, 42, 16, -29, 29, 41, 18, -27, -19, 44, -16, -13, -1, 67, -12, -19, 28, 1, 48, 3, 36, 9, 54, 32, -28, 20, 1, -28, -11, -16, -37, 34, -10, 10, -12, -24, 22, -17, 22, -32, 10, -13, -9, 7, -7, -15, -6, 13, 10, -26, -29, -11, 4, 0, 21, -35, 25, -12, -4, -22, 29, 47, 2, 9, 18, 12, 38, -11, -35, -16, -24, -18, 4, -9, 29, -21, -26, 22, -45, 5, -18, 16, -26, 34, -2, -1, 53, 26, -34, 5, 44, -7, 24, 10, 18, 6, -11, 40, 32, 41, 27, 52, -29, -8, 11, 16, -32, 16, -20, 3, 23, 9, 22, 33, -2, 18, -20, -1, 21, -8, 38, 36, -34, -38, 38, -26, -15, 40, 8, -30, 30, 23, 47, 26, -3, 27, 5, 32, 8, 37, -8, -15, -25, 23, 29, 9, -5, 13, -12, 16, -41, 6, 4, 15, -32, -7, 16, 6, -13, 35, 11, 34, 19, 23, -23, -21, 24, 30, 34},
  '{-27, 8, 26, 26, 4, 20, -29, -2, -1, -11, -31, 15, 17, 33, 17, 22, 40, 5, 27, -15, 4, 16, 28, -6, 8, -11, -21, -26, -32, -33, -27, 4, -26, -55, 25, 35, -4, -31, 50, 0, -20, -12, 6, 17, -36, -9, -7, 26, 29, 24, -27, -2, 25, 16, -10, -19, -2, 29, -17, 14, 1, -9, 11, -17, 4, -38, 5, -18, 40, -10, -4, 24, 26, -15, -32, 4, 2, -5, 24, 14, -7, 18, -34, 41, -23, -5, -15, 14, -21, -65, 8, -35, 36, -28, -20, 15, -28, -20, 1, -5, 38, 25, 27, 1, 34, -7, 8, -5, -3, -10, -3, 8, -10, -24, 0, -5, 11, 6, -32, 14, 0, -14, -3, -8, -32, -20, -13, 33, 46, 23, -16, 1, -44, 18, 19, 6, 7, 43, 42, 54, -19, 2, 26, 21, -15, -7, 12, 15, 3, -11, -25, 21, 3, 34, -31, -10, 2, -7, -4, -8, -2, -36, 37, -9, -16, 15, 5, -7, 9, -10, 35, -40, -11, 30, 1, 25, 6, -4, -16, -7, -10, 17, -28, 30, 22, -10, 21, -24, -8, -38, -5, -24, 17, 25, 10, -2, -7, -42, -7, -9},
  '{9, -8, 8, 31, -21, 0, 26, -21, -12, 24, -13, -4, 11, -16, 4, -6, 1, -3, -25, -21, -21, 29, 13, -4, -12, -39, -22, -28, -17, -24, -65, -1, 2, -34, -22, -83, -40, -53, 29, -61, -40, -85, -49, -54, -47, -38, 37, 17, 14, 25, -29, -9, -18, 22, 13, 29, -10, -38, 1, 12, 44, -22, -7, -5, 27, -9, -14, -21, 1, 20, 34, 33, 36, -46, -34, -14, -14, -12, -4, 2, -23, -26, -9, 39, 6, -14, 33, 30, 19, 55, -18, 41, -16, 44, 48, -19, 5, -24, -38, -29, -2, -36, -29, 18, -5, 31, -15, 35, -31, 4, -8, 36, 3, -28, 50, 8, -20, -30, -7, 47, -30, 34, 28, 36, -37, -8, -4, -15, -31, -27, -29, -32, 11, 15, -16, -2, -35, -31, 28, -25, 1, -39, -8, -17, 29, 11, 30, 29, -20, -15, 0, -23, 29, -4, -24, 11, 34, -11, 27, 32, -14, 37, -35, -14, -1, -9, -19, -32, 16, 41, -16, 8, 36, 43, -21, -30, -12, 20, 33, -4, 14, -35, 5, -32, -14, 54, 10, 14, 0, 28, -20, 37, 7, 2, 7, -5, -29, 8, 9, 14},
  '{0, 4, -7, -13, 10, 2, 0, 5, -8, 15, -3, 0, 20, 3, 0, 7, -4, -6, -5, 4, 17, 7, 3, 4, -2, -2, -4, 0, -4, 0, 0, -2, 0, 2, -11, -1, 0, 9, -4, 6, 0, -1, 4, -3, -1, 1, -2, 0, 0, -9, 0, 2, 0, 1, 4, 0, -6, 0, 7, -3, -2, 0, 0, -9, -7, -12, 0, 0, -2, -1, 7, -13, -3, 4, 0, 0, 6, 12, -9, -3, 0, -2, 12, 1, 0, 0, -14, 0, 1, 0, 11, 0, 0, 1, 1, -10, -10, 0, 8, 0, 1, 6, 12, 8, -1, 1, -12, 9, -3, 16, -11, 0, 1, 11, -11, -17, -1, -6, 3, -3, -7, -20, -5, 0, 20, 0, 1, -1, 12, 0, 0, 2, -6, -1, -18, 0, -1, -2, 1, 0, -1, -5, -16, 3, 0, 5, 8, -10, 11, 1, 0, -9, -9, 18, -1, -1, -2, -12, 12, -4, 5, -1, -3, -5, -9, 12, -1, -1, -1, -16, 12, -1, -18, -3, -4, 1, -13, 12, -18, -13, 1, -5, -10, 7, 2, -1, 7, -4, 22, -15, 8, 10, -18, -14, -6, 0, 8, -20, -18, 13},
  '{21, -3, -11, 37, 27, 28, 0, -11, 16, 38, 7, -27, -5, -16, -8, -28, 7, 19, -28, -34, -12, 18, 41, 32, 10, -10, 13, 20, -5, -31, -1, -26, -43, -12, 0, -47, -15, 34, 38, -22, 24, -23, 11, 15, -5, 14, 5, -34, -34, 35, -10, -23, 34, 21, -42, -1, 20, 9, -19, 30, -1, 26, 33, 31, 3, 16, -11, -6, 23, -13, 14, -47, -19, -46, -13, -11, -11, -20, -9, -1, 4, 0, 18, -4, 11, 5, -11, 3, 25, -3, 26, 27, -28, 22, 31, 1, -43, -13, -13, 18, -40, 7, 22, -26, -27, -46, -10, 23, 16, -4, 12, -28, -6, -36, 41, -24, 11, -49, -19, 14, 25, 25, 23, -41, -9, 33, 5, 30, -12, -8, 10, -19, 6, 28, -12, 23, -18, 9, 36, 9, -11, -3, -28, 23, -5, 31, 15, -36, -25, -24, -41, -39, -40, -33, 1, -28, 26, -25, 15, 4, 6, 18, 25, -23, -2, 19, 16, -44, 2, -3, 2, 19, 15, -13, -26, -42, -6, -31, -30, -18, -27, 7, 36, 34, -5, 26, 37, -21, 3, 13, 42, 32, -2, -13, 32, -24, -33, -26, -18, 3},
  '{-29, 30, 48, 4, 42, 36, 25, -13, 33, 23, -10, 23, 3, -39, -19, -6, 18, 15, 4, 32, 14, -30, -14, -41, -13, 14, 68, 3, -26, -26, 74, 15, 72, 35, -55, 32, 24, 51, 15, 15, 8, 26, 5, -40, 71, -43, -37, -7, -31, 49, 7, -9, -40, -9, -18, -37, 13, 39, 36, -5, 1, -29, 30, 34, -13, 18, -42, -35, -21, -10, -21, 5, 7, -22, 18, -23, -31, -51, -42, -49, -20, 4, 12, -34, -3, -31, 4, -7, -8, 33, -18, -3, 19, 28, -28, -21, 36, 8, -29, -63, 19, 26, 1, 29, -23, 33, -4, 33, -1, 18, 2, 10, -28, 21, -4, 14, 7, -14, -33, -1, 1, -32, 29, 13, -32, 22, 33, 48, 37, -28, 11, 68, 74, 73, 6, 14, 16, -41, -3, -23, -25, -28, 7, 3, -6, 8, 9, -3, 7, 40, -13, 20, -24, -8, 16, 31, -14, 34, -17, -7, -37, 3, -43, -14, 6, 23, 12, -5, 46, -20, 12, 28, 3, -7, -22, 4, 23, -20, 32, 23, 4, -7, 34, -22, -7, 33, -2, -5, 9, 26, 26, 35, -38, 23, -18, 15, 15, -39, 10, -36},
  '{0, -23, 8, 38, -29, 17, 15, 24, 44, 10, 13, 21, -44, -5, 27, -15, -12, 30, 8, 23, -3, -17, -56, 30, -20, 36, -2, 10, -36, 18, 35, 63, 23, -79, -25, 10, 17, 32, 17, -16, 4, 25, 49, 20, -14, 23, 46, 8, 23, -7, 17, -12, 15, 77, 25, -6, 27, 54, 1, -12, 46, -28, 36, 43, -37, 38, 7, -20, 11, -29, 9, -12, 2, 27, 55, -6, -10, -7, 25, 34, 21, 19, 32, 23, 21, -1, -30, 25, 76, -20, -15, 19, 24, 19, 12, -22, -10, 38, 21, 18, 25, -9, -25, -17, -21, 32, 8, 23, 6, 10, -6, -35, -14, -12, -29, 17, -21, 35, 5, -26, -41, -6, 27, 34, -35, -4, 28, 15, -61, -42, -10, 1, -5, -9, -30, -9, -47, -14, 30, -8, 28, 3, 1, 37, 14, 17, -27, 38, 48, -19, -36, -28, -38, 45, 14, 11, -4, 24, -3, 2, 3, -15, 29, 59, -26, 30, -29, -12, 31, -31, 6, 13, -25, -15, -24, 13, -13, 20, 15, -16, -19, -26, 24, 13, 20, 1, -32, 5, 51, 14, 29, -40, 16, 1, -33, -8, 14, 10, 25, 21},
  '{-16, 18, 12, 21, -4, 1, 4, -24, 23, 4, 2, -1, -6, 6, -16, -1, -2, 9, 0, 10, 0, 2, -19, 21, -8, 1, 0, 0, -1, 3, 3, 13, 10, 1, 4, -2, -2, 14, 3, -2, 4, 3, -2, 0, 4, 1, 2, 0, -7, 9, 3, -3, 0, 0, 0, -1, 7, 2, -5, 0, -1, -7, 13, -10, 0, -1, 0, 5, 12, -1, 0, -9, -1, 4, 0, -1, -9, 0, 0, 0, 0, -10, -2, -2, 0, 0, -1, -2, 10, 0, 0, 0, 2, 5, 0, 0, -3, -2, -9, 0, 10, -22, -13, -13, 1, -12, 19, -20, -17, 8, -2, -2, 5, 0, -7, 0, 0, -17, 1, -18, 0, 1, 19, -13, -3, -1, -1, 0, 0, 0, 2, 14, 6, -10, 0, 0, -5, 3, 11, 5, 0, 0, -6, 2, -1, 0, 0, -1, -10, -7, 1, 18, -1, -1, -2, -3, 9, -11, 23, -11, -1, -1, -15, -1, 13, -1, 0, -18, 26, -14, 0, 2, 12, -6, -11, 11, -11, -16, -19, -4, 2, 6, 21, 13, -4, -2, -2, -24, -25, -21, 0, 0, -11, -21, -19, 0, -1, 0, -15, -18},
  '{9, -7, 47, -14, 12, 30, 2, -11, 43, 5, 26, -17, -34, -46, -29, 8, 46, 23, -9, -2, 18, 33, -53, -23, -30, 6, -21, 20, 9, -37, -16, 50, 22, -19, -33, -4, 32, 37, -2, 12, -7, 23, 56, -27, 7, 13, 18, 18, -16, -41, -11, -37, -5, -32, -21, 1, 4, 22, 18, -5, 20, 16, 0, 59, -12, -31, 31, 38, 31, -40, -4, 23, -5, 3, -9, -33, -10, -3, -6, -29, 12, 4, -27, 8, -12, -37, 19, -23, 3, -2, -22, 16, -8, 65, 2, 14, 13, 44, 32, 1, -27, -39, 16, -20, 26, -30, 36, -1, 59, -16, 2, 19, -30, 2, 6, -14, -40, -53, 31, -24, 32, -7, -9, 18, 11, -1, -32, -7, -52, -38, 28, 11, 58, 42, 22, -23, 17, 34, 26, -30, 56, 15, 31, 36, 12, -1, -53, -10, 9, -12, 32, 20, 27, -32, 26, -11, 37, 38, -1, 38, -22, -2, -11, -37, -21, -32, 21, -21, -9, 3, 27, -23, 23, -3, -47, -16, 10, -10, 15, 4, -15, -10, 22, 35, 13, 6, 19, -18, 13, 21, 33, -8, -34, -20, 33, -25, 0, 14, -37, -45},
  '{9, 1, -3, 19, 3, 20, -10, -28, 1, -21, 8, -8, 40, 64, 54, -5, -5, 20, -44, 13, -18, 34, -21, 16, 55, 12, 41, 32, 24, 90, -45, -15, 40, 60, 38, 36, 0, 27, 51, 48, -25, 5, 56, 2, -25, 38, 8, 8, 46, -11, 33, -20, -26, -29, -30, 38, -15, 19, 11, 17, 38, 17, -9, -12, -15, -21, -24, -3, -8, -11, 12, 13, -42, 30, 6, -13, -26, -13, -42, -60, 11, 25, -35, -31, -36, 35, -23, 12, -24, -28, -18, -43, -42, -38, -6, 17, -15, -18, -8, -4, -13, 20, 50, -16, 10, 0, -11, 18, -26, 22, -31, 2, 4, 16, -20, 17, 12, 41, 20, 33, -23, 16, 31, 27, 16, 8, 8, 32, 25, 54, -19, 48, 31, 36, 34, 8, 1, -2, -19, 22, 8, 41, 8, 33, -19, 26, -11, 32, -14, 11, 2, 21, -20, 42, 19, -22, 25, 34, 20, 7, 11, 19, -29, 2, -14, 19, 21, 42, -15, -30, 45, -10, 28, 14, -11, 8, -14, 33, -13, -25, -12, 5, -17, -36, -21, -32, -9, 19, 6, -6, 5, 1, 38, -20, -24, 37, -20, 20, -22, 50},
  '{-18, -13, 35, -39, -32, 5, -1, -30, 0, 27, -16, 9, 13, -10, 20, -14, 7, 2, 42, -16, 46, 34, 66, -18, 10, -32, -13, 25, -14, 30, -10, 31, 9, 13, 5, -7, -35, -22, 59, -26, -7, 28, 40, 25, -47, 18, 1, 13, 53, 25, -7, -28, -33, -39, 8, -27, 5, 13, -15, 1, -31, 24, -8, 21, 15, -19, 1, -4, 9, -2, -37, -24, 11, -41, 11, 20, -22, -17, 15, 4, 16, -23, -27, -8, -34, 6, -13, 40, 9, -27, 4, 30, -47, -33, 32, -14, 14, -15, -1, -2, 41, 36, 0, 10, 24, -3, -45, 2, 40, -45, -44, 18, 10, -52, 25, -33, -7, -47, 14, 45, 40, 11, 30, 20, 46, 10, 17, 47, -29, -26, 14, -19, -8, -12, 39, 7, -23, -10, 5, 9, -42, 36, 4, -46, -12, 7, -1, -9, -5, 21, -8, 30, 10, 25, -39, -13, 15, -23, 39, -29, 27, 39, -8, 7, 9, -19, 12, 11, -3, 25, 3, 9, 44, 12, -15, 6, 34, -3, -27, 27, -8, -42, 7, 36, -24, 1, 0, 7, -25, 14, 17, 8, -29, -12, 17, -7, -15, -15, -6, 7},
  '{31, 30, -16, -2, -40, 18, 34, 10, 24, 31, -9, 32, -36, 14, 30, 5, -8, 9, 6, 17, 46, 22, -11, -43, 3, -22, 37, 28, 11, -11, 19, 13, 16, -10, -31, -7, 8, 1, -17, -39, 32, -3, 20, -25, -12, -32, 9, 17, 10, 44, -6, -18, -6, 19, 21, 24, -5, -3, -3, -12, -18, -5, 28, 17, -37, 3, 15, -38, -6, 7, -9, 13, 17, -3, -34, -27, 23, 20, 15, -16, 3, 6, 21, 7, -11, -28, 9, 2, 15, 28, 17, 0, 20, -2, 47, 7, -12, 24, 1, -18, -3, -9, -19, 30, 0, 2, -3, -28, 25, 5, 25, 10, 0, -30, -2, 21, -39, 27, -37, 0, 3, 6, 17, -34, -26, 29, 23, 2, -43, 5, 7, 35, 24, -25, -40, 9, -25, 18, 25, -22, 38, -14, -17, -22, 6, -26, 19, 26, 2, -15, -18, 5, -33, 40, -23, -7, -19, -20, 49, 29, 5, -35, 25, 13, 0, 15, -20, -11, 20, 47, 9, 0, 19, 12, -36, 22, -21, -9, 23, -6, 7, 15, 31, 29, 3, -25, -6, 3, 6, -16, -30, -28, -17, -3, -21, 24, -37, 21, 0, -31},
  '{43, -37, 17, -45, 4, -20, -21, -17, 38, 19, 7, 42, -52, -44, 28, 9, 31, 25, 39, 51, 61, 14, 26, -27, 4, -25, 33, 40, 46, 6, 45, 59, 36, -45, 3, 16, 10, 11, 39, -60, 31, 53, -6, -7, 8, 32, -8, 74, 23, -8, 6, 0, 14, 51, 44, 6, 19, -7, -33, -36, -14, 0, 1, 25, -34, 17, -30, 19, -38, 23, 11, -2, 13, -11, 4, -22, 26, 21, 37, 45, 14, -27, -3, 72, 13, -33, 3, 3, 55, -42, -7, 20, 28, -11, -35, 18, -12, 33, -42, -49, -10, 2, 16, -7, 16, 12, 1, -20, 5, -33, -40, -42, 9, -14, 2, -29, -2, -21, 29, 18, -20, -34, 3, 11, 10, 47, 64, -11, -16, -19, 8, 21, -11, 2, 2, -17, -45, -37, 5, -27, 6, -22, -19, -31, 48, -27, 7, 25, 27, -20, 35, -33, -18, 27, -28, 12, -11, 10, 11, -28, 6, -31, 24, -17, -44, -25, -11, -30, -14, 26, 33, 17, 44, -26, -28, 12, 18, -39, 30, 15, 0, -23, -24, 42, -30, -7, -17, 34, 34, 32, 18, 21, 40, 20, 45, 19, -34, -20, 8, -27},
  '{19, 26, 1, -32, 7, 12, -29, 3, 2, -3, 13, -23, -24, 15, -28, 30, 15, -9, -7, 17, 34, -35, -16, -2, -33, -9, -37, -8, -14, 2, 26, 20, 49, -22, -8, 38, 64, 5, -21, 0, 20, 41, 3, 43, 52, -26, -35, -38, -44, 40, 13, -3, 14, 14, 24, -19, -17, 12, 35, -24, -31, 30, 48, 38, 7, 36, -8, -24, -40, -14, 17, 15, 37, 39, 1, 19, -20, 6, 23, 46, 7, 12, 17, 9, 46, -29, -14, -7, 0, -5, -9, -16, 6, 17, -44, 28, 0, 14, 12, 6, -12, -14, -15, 2, -16, -29, -33, 17, -21, -3, 21, -16, 18, -14, 25, 5, 17, 27, 19, 20, 13, 3, 34, 0, -4, -3, 60, 47, 21, -16, 53, 19, -8, -1, -20, -11, 18, 4, 19, -33, 19, -36, -28, 15, 54, 26, 25, -16, -31, -28, 22, -16, -14, -26, -25, 9, -41, 18, 33, 17, -11, 20, 28, 20, -8, 21, -14, 38, -33, 8, 28, 32, 20, -11, -50, -24, 41, 9, -8, 10, -40, -43, 22, -1, -30, 4, 12, 17, 9, -28, -9, -36, 25, 34, -39, 45, -18, 14, -26, -50},
  '{11, 2, 46, -22, 3, -10, 29, 13, 23, 1, 13, -3, 5, 21, -12, 61, 18, -12, 7, 39, 8, 2, 36, 41, 32, 30, 14, 2, 14, -47, 62, 46, 86, 7, -51, 67, 72, 30, 5, 72, 34, -7, 28, 1, 2, -8, -19, -9, 19, 4, 24, 11, -35, -11, 30, 4, -10, 31, 27, 1, 18, 16, -2, 24, -24, -4, -4, -21, -45, 14, -9, -60, 10, 0, 7, -2, -5, -44, -42, -4, -9, 10, -39, -23, 20, -7, -31, 13, -10, -42, 14, 21, 7, 2, 5, 16, -38, 11, -29, 9, -19, 13, 14, 13, 27, 33, -22, 1, 37, 45, -31, -31, 20, -13, 16, -8, -16, -34, 27, 16, 21, -10, -31, 9, 42, 10, 17, 5, 5, -7, 28, 10, 78, -2, 39, -17, 15, 20, 3, 0, 23, -9, 28, -16, -10, 30, -10, 4, -10, 26, -25, -1, 0, 34, -4, 24, -37, 31, 44, -3, -25, -17, -5, -11, 1, 13, 16, -4, -37, 24, 44, 24, 34, -6, 33, -14, 30, -14, 43, -22, 32, -12, -14, 26, -14, 4, -37, -13, -4, -20, 26, -15, 33, 2, -11, 27, -8, -29, -20, -8},
  '{18, 17, -23, 18, -35, 46, -35, -30, 5, 13, -31, 22, 18, 28, -13, -19, 2, 3, -19, -6, -47, -26, 0, 47, -16, -13, 12, 21, -34, -26, 30, -1, -16, -13, 1, 34, -27, -17, -42, -41, -30, -30, 18, -41, 10, -46, -21, -12, 15, 41, 2, -17, 24, 0, 32, -33, -18, 42, -29, -13, 6, -13, 5, -62, -39, -23, 22, -8, 23, 13, -45, -22, -17, 28, -20, -18, 25, -14, 10, 7, 10, 19, -10, 6, -1, 16, -29, -18, 12, 36, 32, 27, 32, -51, 23, -21, -8, -5, -30, -10, -28, -15, -5, 56, -16, -22, -4, 33, 10, -43, -35, -12, -20, 34, 33, 9, 11, -19, 43, 2, 2, -24, 24, 27, 34, 20, 35, -22, -2, -14, -32, 10, -35, -19, -4, 35, -14, -15, 25, 22, -14, -19, 17, -21, -34, 15, -29, 23, -16, 25, 0, -32, -3, -4, -32, 31, -9, -17, -26, -37, -17, -37, 47, 53, 7, 22, 26, 28, -19, -15, -9, 22, -1, 19, 4, 22, -20, 32, -20, 21, 3, 2, 35, 33, -31, 0, 2, 20, 52, 11, 11, 38, 54, 8, 32, -39, -24, -16, 29, 41},
  '{-2, 1, -1, -1, -2, 2, 0, -2, -2, -4, -1, -2, 0, -7, -6, -4, 0, 1, 19, 1, -1, -1, -11, -7, 11, -1, 0, -2, -2, 1, -1, 1, -4, 0, -2, 0, -5, -1, -1, 0, -4, -7, 0, 0, -1, -1, -1, 2, 1, -1, 1, 0, -9, 1, 1, 0, 0, -8, 0, -3, 0, 0, 0, 0, -3, 0, -2, 6, 0, -3, -3, -4, -12, 1, -1, 1, 0, -1, 0, 1, 8, 1, -7, 0, -1, 0, 0, -8, -1, -2, -1, 0, 1, -2, -1, -2, -4, 5, -1, 2, 0, -11, -9, -18, 0, 0, -1, -21, -3, -1, -1, -1, 5, 4, -1, -1, 0, 15, -1, -5, -1, -8, 6, -7, -9, -1, -1, -1, -1, 1, -2, 0, -5, 13, 0, -1, 17, -6, -3, 0, -2, 0, -14, -2, -1, -2, -5, 10, -2, -5, -1, 9, 16, 3, -1, -15, 17, -14, -1, -6, 13, -6, 10, 14, -1, 3, 0, -12, -4, 2, -2, -1, 20, -1, 1, 1, 9, 4, 13, 3, 8, -1, -1, -1, 1, 3, -1, 4, -1, -9, -2, 0, -17, -1, 0, -2, -9, -10, -5, -4},
  '{-20, -25, 25, -30, -3, 13, -8, -47, 7, -7, 25, -39, 18, -11, 35, -11, 20, -20, 9, -30, 20, -4, 1, 31, -32, -31, -15, -20, -26, 6, 8, 0, -40, -15, -32, -17, -38, 9, -14, -14, 26, 33, -15, 5, -44, -19, 28, -2, 11, -31, 30, -16, 19, 25, 7, -19, -17, 11, 24, -33, 39, -19, 5, -19, -17, 14, -5, 44, -6, -10, -20, -30, 5, 26, -11, 0, 25, 42, 46, 13, -13, 39, 33, 37, 3, 1, 8, 31, 22, 11, 2, -18, 30, -24, 22, 2, -17, 15, 5, -4, -3, 29, -26, -4, -10, 37, 32, -21, 10, 14, -3, 17, -25, 32, 0, -5, -18, 10, 12, 16, -21, -29, -13, -31, -32, -3, 15, -38, -27, 27, -11, -7, -19, -6, -26, 16, -2, -4, 21, 29, 14, 38, 43, 16, 6, 0, 16, -26, 40, -40, -20, 18, 9, 17, 31, -7, 12, -34, 18, 11, 7, -4, 8, 43, -20, -2, 22, -9, -1, 37, 17, 18, 10, 33, 0, 20, -15, -28, 0, 33, -23, 8, -6, 4, 22, 27, -11, -14, 0, 3, -24, 21, -14, 6, 27, -33, -4, -21, -14, 27},
  '{27, 14, 6, 22, -38, 15, -13, -50, 15, 15, 24, -26, -23, 27, 24, -20, -1, 19, -5, 31, 3, -1, -10, -27, -27, 13, -20, 32, 5, 53, -33, 3, 31, -44, -34, 10, -42, 10, 20, -17, -22, 34, 51, -14, -47, 43, 48, 29, -16, -12, -37, -25, 13, 10, 17, 27, 16, 29, -1, -33, 24, -39, -41, 11, 2, 25, 29, 25, 31, 34, 24, 35, 9, 30, 6, -5, -3, 0, 24, -21, 10, 23, -26, -29, -1, -12, -4, 2, -16, -49, 22, -28, 11, -4, -19, -1, 8, -30, 22, 13, 38, 18, -29, -17, -18, -8, 8, 20, -36, -41, -23, 39, -1, -9, -25, -17, -16, -15, 23, 16, 29, 8, 10, -1, 4, -30, -6, -6, 2, 7, 23, -16, -4, 7, 9, 17, -5, -12, -21, -8, 5, -8, -19, 15, -3, 3, -8, -24, 29, -2, 40, -18, -16, -2, 2, -9, 3, -19, -7, -5, -5, 30, 21, -20, 50, -38, -25, -26, 14, -14, -33, 24, 14, 31, 8, 39, -13, -11, 35, -6, 0, -22, 13, 7, 31, 25, -1, 14, 25, 52, -36, -16, 9, -4, 49, 1, 34, -38, 3, -17},
  '{-39, -17, 4, 25, -31, 22, 0, 25, 3, 49, 28, 25, -15, 5, 34, 23, -12, -10, 24, 18, 13, -4, 14, 14, -66, -40, -1, -26, 23, 65, -14, 46, -9, 48, 59, -18, -67, -20, 5, 30, 5, 1, -27, -50, -12, 17, 4, -30, 37, -24, -24, -7, 10, -9, -10, -12, -7, -26, -18, 35, 8, 10, -7, -27, 27, 8, 26, -23, -4, 43, -14, 33, -32, -4, -39, 25, 8, 12, 7, 8, 8, -28, 9, -34, -48, 10, 2, -5, -21, -26, -6, 12, 3, -10, 14, -12, 33, -28, 15, -15, 46, 2, 14, 1, -30, 17, 19, 16, 28, 1, -25, 46, -10, -26, 27, 23, 22, 25, 8, 8, 27, 43, 3, -22, 17, -23, -5, 23, 46, 17, 3, 15, 23, 53, 56, 10, -17, -11, -16, 40, -5, 25, -1, -41, -26, -17, -11, 27, -25, 0, -22, -20, 17, 6, 28, -31, 30, -4, 31, -17, 29, -26, -10, -35, 34, -8, 7, 19, 14, -1, -15, -10, 18, 17, -30, 2, 35, 30, -30, -17, 34, 41, 13, -3, -20, 18, -6, 3, -5, 13, -8, 40, -28, -40, 25, -36, -13, 37, -22, 9},
  '{-13, 16, 51, 30, 29, 28, -6, 22, 8, 23, -36, -9, 41, 37, 46, 26, 8, 31, 8, -10, 3, 5, 8, 1, -47, -3, -19, 11, 42, 26, -27, -11, -18, 8, 43, 18, 18, 47, -8, 33, 71, 40, -4, 29, 5, -10, -30, -50, -48, -40, 9, -28, 9, -30, -28, 34, 44, -34, -8, -4, 18, 27, -1, 1, -3, -7, -12, 48, 56, -19, -20, 12, 38, 11, -11, -5, -21, -9, -58, -12, 2, 29, -2, -60, 36, 14, 1, 5, -15, -51, 39, -23, -24, 53, -17, -17, -40, -9, 39, 42, 34, 16, 23, -29, 13, -18, 49, 40, -17, 41, -22, -3, 12, 11, 20, 27, -33, -23, -16, -32, -34, -11, -35, 15, -50, -18, -50, -9, -11, -9, 9, 3, 15, 32, 16, 34, 33, 55, -7, 23, 50, 28, 27, -2, 20, 2, -3, -7, -6, -12, -33, 24, -17, -14, 34, 8, -3, -22, 11, -15, -31, -34, -26, 4, 17, -39, -9, -17, 16, 15, -28, -8, 35, -8, 5, 45, 26, -8, -27, 31, 5, -9, 10, 0, 46, 38, 26, 8, 25, 45, 14, 0, 18, -32, 23, 30, -20, -8, 14, -5},
  '{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
  '{-2, 42, -11, -15, 7, -37, 13, -9, 18, 0, 36, -33, 22, -12, 29, 1, 29, -16, -1, 27, 25, -11, 63, 38, -16, 3, -31, -23, 1, 30, 3, 21, -2, 21, 7, 26, 2, 20, 44, 59, 4, -27, 8, -26, -28, -31, -3, -2, -36, 18, 40, 31, -45, -38, -67, -31, -18, -26, -3, -11, -9, -15, -3, 5, 60, 8, 31, 17, 26, 17, -33, 27, -15, -14, -26, -5, -2, -6, -24, -17, -33, -10, -27, -34, 7, 7, 20, -2, -51, -15, -39, 52, -33, 3, -30, 1, 32, -5, -8, -33, 33, 20, 1, 13, 23, 15, 40, -17, 10, 26, 20, 41, 4, 15, -8, 6, 17, 18, 10, 10, 32, -6, 29, 21, -6, -26, -22, 9, -5, -37, 38, 25, 27, 10, 58, -14, -17, 30, 24, 36, -14, -33, -17, -26, 23, 29, 38, 22, -4, 12, 32, -26, 45, 14, -21, 26, 10, -11, 4, -14, 19, -18, -38, -33, -11, 25, 33, -3, -22, 49, 29, -15, 12, 30, 6, 9, -27, 0, 21, 7, 40, 43, -3, 7, 6, -22, -15, 10, -51, 15, 34, 12, -16, -38, 36, -35, -5, 26, -20, 29},
  '{7, 23, -10, 13, -3, 6, -10, -23, -9, -24, 25, 8, 27, -4, -12, -9, -11, 12, -3, -16, 0, 1, 0, -3, 14, -7, -3, 8, -8, 6, -2, -1, -9, -3, 0, 0, 3, 3, -1, 0, 13, 16, -2, 2, -2, -16, 6, 1, 7, 4, -4, -1, 0, 1, -8, 1, 0, -1, 9, -7, -16, -1, 0, -10, -4, 6, -9, 1, 6, 0, -4, -3, -2, -7, -9, 0, 0, 0, -1, 1, -1, 0, 0, -1, 6, -1, 0, 0, -1, 0, 2, 0, 0, -1, 0, 0, 0, 0, 5, 0, 0, -15, 1, -16, 17, -15, 24, 4, 10, 6, 26, 6, -25, -11, -25, 24, -12, -30, 16, 24, -6, -7, -7, -24, -9, 0, 0, 0, 0, 0, 4, -1, 0, -2, 7, -15, 8, -2, -1, -8, 12, 18, -2, -12, 2, 4, 0, 2, -7, -5, -1, -18, -5, -12, 1, 4, -5, 3, -7, 6, -20, -21, -16, 11, 0, -9, 17, 21, -16, 12, -1, 0, 0, 5, 3, -4, 15, -2, 7, -23, -6, -27, 19, 7, 2, 24, 2, 9, -26, -18, 6, 7, 10, -16, -1, -3, -11, 4, -8, 0},
  '{-34, -7, -14, -32, -14, 6, -26, -14, 0, 49, -6, -24, -16, -35, 33, -34, 34, 14, 14, 46, -8, -36, 63, 35, 4, -34, -37, 2, -6, 13, -55, -20, -62, 24, 20, -31, -58, -44, 7, 22, 6, -73, -6, -38, 19, -20, -55, -56, -32, -9, -22, 10, -29, 8, 20, 37, -7, -42, -42, 7, -26, 22, -21, -17, 34, -10, 17, -7, -19, -16, 25, 1, -6, -43, -22, -13, 28, -10, -8, 29, -24, 32, -22, -23, 15, 1, 41, -7, 11, -3, 10, 32, 7, -10, 15, 28, 29, -6, -10, 0, -6, 18, 27, 31, 40, -1, 18, 11, -23, 2, 33, 42, 21, 5, 48, 8, 21, -2, -17, 12, 6, -12, 14, 38, 37, 25, -30, -13, 2, 55, -24, -10, -52, -4, 9, 8, 31, 19, -17, 45, 7, -15, -29, -44, 19, -23, -16, 10, 31, 29, 1, 0, 34, 18, -14, -12, 42, 18, 28, -19, -18, -7, 29, -16, -14, 34, 39, 15, 7, -21, 5, 14, -1, 31, 2, 6, 10, 0, 14, -19, 2, 38, 3, -24, -6, 22, -10, 2, -42, -7, 10, 0, -15, -26, -19, 15, 12, -13, -9, -33},
  '{3, 16, -9, -16, -21, 20, 26, -21, 1, 2, 15, -10, 20, -13, -29, 38, -9, 16, 13, 0, -13, 3, 8, -36, 27, -15, 56, 8, -53, -75, 64, 43, 11, -45, -85, 8, 72, 4, -18, 14, -24, 70, 38, 26, 16, 47, 25, 26, 26, -17, -16, -39, -11, 55, -9, 21, -9, 8, 14, -4, 15, 20, 30, 21, -15, -38, 22, 49, -22, 15, 9, 6, 1, -14, 3, 0, 5, -4, -34, -45, -34, -21, -25, 18, 12, -13, -16, -43, 46, -10, 8, 5, 9, -6, 2, -18, 9, 37, -28, -24, 30, 25, 32, -18, -12, 3, 24, -19, 32, 26, -2, 8, -4, 17, 33, -31, -23, -10, 15, 0, 8, -1, -13, 10, -3, -18, 17, -7, 28, -29, 47, 30, 24, 5, -58, 0, 11, 31, -34, -44, -28, 2, 60, 15, 35, 26, -9, 3, -26, 18, -17, 17, 12, -6, 18, 16, -4, 24, 48, -19, -33, 2, 43, 0, 40, 1, 16, -16, -15, 15, 21, -24, 6, -5, 8, 4, 22, -26, -21, -3, 8, 35, -8, 27, -5, -13, 23, 13, -5, -20, -12, -22, -3, 14, -20, 32, 3, -38, -9, 34},
  '{31, 17, 15, 61, 29, 44, 38, 55, 58, 12, -10, -10, -41, 10, 8, -41, 50, 27, -32, -24, -2, -35, 24, -46, -28, 25, 28, -4, -21, 1, 19, 4, 55, 24, -54, -21, -4, 18, 16, -27, -48, -41, 21, -42, 4, 2, 19, -32, 27, 44, -40, -8, -46, -40, -37, 3, -16, 3, -5, 27, 26, -37, 21, 43, 60, 19, 31, -50, 19, -11, -25, -5, -28, -6, -6, -17, -23, 12, -33, -58, -36, -18, -15, -34, -48, 8, 10, 35, -17, 27, 6, 5, -4, 5, 31, -4, 25, 11, -11, -32, 22, 33, -10, 7, -3, 33, 39, 39, 9, 18, -20, 29, 14, -9, 33, -31, 9, -5, -36, 31, 17, -5, 10, 15, 12, -20, -20, -33, -19, -16, -27, -14, -5, 14, 24, 2, -6, -27, -8, 24, -22, 7, -36, -19, 10, -36, -26, -13, 12, -30, -11, 30, 34, -10, -13, -16, 17, 8, 53, -15, -20, 3, -42, 17, 22, 37, 32, -26, -30, -22, -38, -26, -20, 34, -51, -41, 21, -16, 27, 32, 29, 41, 32, 19, 51, 27, -25, -10, 0, 53, -6, -25, -19, 2, 12, 31, -15, -11, 11, -42} 
};

reg  signed [7:0] fc2_weights_re[10][64] = '{
  '{40, -8, 35, -60, -23, 24, 76, 67, -97, 54, 1, -19, -49, -56, 5, -17, -19, 11, 53, -79, -2, 17, -1, -27, 43, 21, -5, 28, 28, 25, 60, 31, 20, -6, 60, -72, 32, -91, -91, 95, 13, 9, 5, -37, 0, 46, -88, 75, 33, 16, -17, -30, -21, 0, -66, -41, 73, -14, 0, 62, 0, 57, -72, 68},
  '{-86, -89, -37, 81, -2, 43, 19, -82, -22, 96, 2, 61, 59, 37, -8, 11, -42, 23, -95, -27, -68, -56, 5, 50, -62, -78, 57, 32, -36, -49, -19, 0, 53, 50, 6, 0, -51, 16, -34, -63, 0, -6, -96, 70, 0, -19, -48, -24, 13, 43, 20, 18, 49, 0, 3, -68, -100, -60, 0, -91, 0, -85, -28, -77},
  '{84, 65, -75, -26, -113, -45, 72, -2, -4, 42, 1, -16, -35, 6, -75, -1, -78, 66, -40, 6, -40, -34, -44, 50, -44, 40, -26, 81, -9, 84, -15, -2, 51, 16, 46, -75, -23, 51, -72, -63, 1, -90, 55, -6, 0, -30, 37, -22, -59, 19, -5, 76, 30, -3, -72, -46, -29, -76, 0, -15, 0, -36, 48, -29},
  '{33, -30, 23, -34, 41, 11, -21, -7, 9, 24, -3, -64, -77, -63, 72, 74, -12, -22, -15, -26, 98, -100, 3, -44, 26, 11, 25, -77, -34, -36, -52, 0, 14, 19, -80, -37, -42, 1, 65, 27, -1, -17, -20, 0, -2, 20, -12, 74, 59, 53, -31, 33, 36, -2, 24, 56, 26, 29, 0, -11, 0, -67, 33, 26},
  '{-19, 74, -60, -41, -43, 35, -101, 79, 57, -14, -3, 53, 78, -26, -98, -27, 84, -9, 64, -66, -108, 60, -77, -83, 68, 29, -70, -39, 6, 8, -11, -7, 49, 85, -56, -58, 57, -41, 28, -13, -1, -123, -78, 22, 1, 24, -75, -68, -56, 29, 0, -88, -13, 1, 72, 12, -50, 52, 0, -56, -23, -1, 27, -96},
  '{-16, 10, 22, 65, 67, 75, 23, 56, 13, -74, -20, 60, -7, 23, 67, -14, -64, 28, -21, -86, -38, 18, 21, -62, -32, 28, 45, -70, 77, -42, -97, 1, -26, -46, -51, -2, 67, -44, -7, -48, 13, -53, -39, -23, 0, 31, 23, 28, -54, 21, -9, -5, -94, -2, -63, -15, 44, 77, 0, 27, 0, -1, -50, -57},
  '{-14, -75, 36, 60, -44, -88, 53, 75, -14, -46, -3, -30, 43, -20, 27, -74, 53, 86, -38, -67, -38, -2, -13, -95, -57, 13, 70, -49, 62, -77, 30, 0, -83, 5, 72, -21, 1, 15, 30, 68, 0, -67, -84, -30, 0, -111, 23, 46, -2, 30, -103, -88, 78, -1, 62, 47, 84, -42, 1, -18, 0, 36, -68, 38},
  '{-53, 19, -3, 36, -18, 29, 34, -7, 24, 73, 4, -35, 66, -78, 81, -90, 0, -81, -51, 67, -84, -64, 36, 71, 22, -79, -96, -39, 4, 63, 1, -59, -70, -16, 26, -104, 19, 21, -45, 3, 0, 16, 84, 35, -12, 61, -63, -47, 20, 63, 46, 50, -31, -8, -29, -41, 23, 72, 0, 7, 2, -11, 0, 86},
  '{66, 41, -66, -15, -75, -15, 31, -31, -48, 38, -15, -33, 64, 42, -73, 49, 43, -15, -31, 19, 15, -14, -16, 50, 59, -70, 73, 73, -90, -67, 29, -1, -83, 67, -84, 1, 13, -18, 37, -26, 0, 45, -20, -54, -1, -73, -19, -91, -87, -94, -3, 9, 51, 5, -48, -55, -13, 81, 0, 26, -1, 27, -17, 14},
  '{33, 53, -98, 81, 58, 69, -9, -11, 43, -10, -2, -1, -30, -18, -77, -73, 24, -101, 36, 71, -25, -31, 9, -28, -18, 70, -43, 18, -28, -9, 81, -3, -33, -57, -25, 46, -25, -48, -41, 15, 0, -83, -17, 32, 0, 62, 37, -49, -19, -71, -85, -75, 60, -5, 57, 27, -37, 38, 0, -70, 1, -110, 28, 77} 
};
*/
reg  signed [8:0] fc1_weights_re[0:12799] = {

-27, -10, -25, -33, 7, -3, -6, 3, 42, 46, 9, 30, 49, 35, 11, 21, 41, 18, -1, -22, 29, 3, -27, -21, -8, 43, -34, -74, -21, -20, 9, 5, -24, -35, -36, 27, -27, 0, 61, 27, 56, -16, -47, 13, 0, 48, 35, -44, 12, 21, -23, 7, -10, -19, -22, -4, -4, -29, -4, -1, 12, 9, -1, 44, 30, -16, 57, -21, -29, 26, 36, 29, -32, -14, -37, -19, -37, -21, 21, -68, 14, 7, 24, -9, 6, -11, 7, 0, 11, 21, 20, 9, -37, 11, -21, 41, -6, -16, -17, 25, 24, -19, -17, -20, -36, -21, 36, 13, 60, 18, 43, 9, -13, -30, 3, -7, -59, -21, 25, -20, -29, -6, 47, -61, -29, 48, 28, 2, -26, -22, -20, 29, -31, -8, 25, -23, -21, 35, 47, 8, 18, -8, -7, 34, 15, 4, 11, -25, -23, -9, -2, 16, -61, 12, -42, -2, -36, -27, -19, 55, 4, -30, 31, 28, 4, 12, 18, 29, -8, -12, -5, 9, -40, -14, -35, 20, 13, -41, -26, -13, -1, 1, 7, -7, -8, 28, -11, 27, 33, 33, 43, 4, -2, -5, 3, -17, 20, 11, -49, 5, 21, -35, 9, 41, 22, -48, -7, 19, 9, -10, -4, -42, 4, 21, -18, -27, 28, 48, -27, 28, 33, 12, 5, -26, 7, 53, -14, 0, -43, 16, -49, -6, 11, -7, 8, -39, -57, -36, -13, -1, -1, -7, -2, -4, -19, -28, 1, 1, 15, 36, -49, 15, -4, 9, 18, -36, -53, 3, -19, -19, -15, -2, 26, 26, -6, 7, 42, -9, -36, -14, 2, -3, -16, -33, -57, -20, 18, 47, 38, 27, 3, -16, 38, 10, -31, -29, -34, -53, -43, 16, -26, 27, 7, 13, 32, 15, -19, 35, -34, 19, 20, 7, 4, -15, 9, -4, -21, -26, -7, -18, 33, 84, -17, 59, -27, -10, -3, -56, -2, 33, -56, -45, 1, 23, -14, 55, 36, 17, -12, 49, 57, 60, 51, -7, -3, -43, -39, 4, 14, -15, 20, 16, 58, 6, 17, -4, -8, -6, -12, 6, 5, 34, 16, 14, -31, -24, 4, 9, 25, -11, 13, -4, 12, 0, 24, 16, 49, 52, -22, 12, 25, 5, 3, -48, 13, -17, 42, 3, 46, -9, -14, -22, 4, -11, 0, 19, -33, -44, -31, 8, -15, 27, -11, 14, 26, -6, 22, 0, -56, -10, -4, -12, -4, 0, 3, 3, -3, 18, 2, -2, 7, -13, 1, 6, -17, 8, 17, 9, -11, -22, 21, 4, -5, -2, 10, -8, -12, 0, -12, 14, -6, -6, 18, -26, 20, 14, -10, 7, -17, 25, 3, -12, 10, -9, 11, -5, -1, 20, 16, -9, -4, -3, 2, 15, 16, 13, 13, 10, -6, -6, 6, -8, -4, -8, -26, 16, 16, 10, 1, 8, 22, -2, -1, 6, 27, -7, -13, -1, -3, 2, -5, -12, 11, 0, 18, -7, -10, 19, -6, -13, 12, -3, -16, -5, -25, 13, -2, 13, 13, -5, 2, 9, 8, 23, 7, 30, 24, 4, -16, -11, -14, -3, -22, -17, -53, 21, 14, 4, 8, 25, 17, -4, -4, 36, 9, -14, -35, -37, -18, 3, -9, -4, 10, 8, 36, -4, -8, -1, -4, -1, -4, -18, -8, -30, -42, 9, 10, 9, -4, 11, -11, 0, -1, -2, 8, 9, 4, 19, 16, -2, 7, -15, -7, -6, -29, 12, 3, -2, -19, 6, 7, -4, -8, 4, 35, -5, -8, -3, 4, 1, 6, 1, 3, -3, 2, 0, 8, 14, -11, -29, 12, 9, -14, -22, -31, 6, 2, -5, 3, 5, -3, -33, 37, -13, -19, 31, -41, -4, 10, -13, -26, 15, 18, -10, -6, 6, -14, 6, -31, -7, 21, 20, -6, 38, 7, -11, -32, -9, -17, -62, -16, -47, -33, 1, -17, -9, -11, 12, -26, 60, 18, 7, -34, 5, 58, -2, -5, 34, -18, -22, -27, -16, 13, -23, 6, 1, 26, 27, 22, -4, 48, -10, 35, -43, -49, -27, 1, 27, 13, -9, -10, -54, 4, 41, 16, -4, -8, -31, 26, 39, -16, 2, 18, 2, 39, -33, -36, -20, -19, -17, 13, -1, 26, 19, 21, -8, -4, 31, 10, -26, -30, 13, 0, 16, -4, 6, 21, 8, -8, 14, -7, 11, 27, 6, 18, -32, 63, 9, -18, -43, 7, 37, 9, -3, -36, -42, 14, -12, 48, 12, -47, -32, -26, 18, 29, -28, -52, -15, 24, 3, -10, 24, 0, 7, -29, -7, 51, 30, 20, -1, 10, 21, 16, 11, -1, 31, -23, 30, -17, -23, 10, -23, 20, 26, 12, 1, 16, -8, -37, -51, -18, 15, 5, 19, 34, 14, -33, 23, -14, 39, -9, 4, 17, -7, -2, -30, 18, 38, 33, 36, 1, 15, -20, 20, 35, -29, 24, 13, -27, 16, -37, 32, -6, 34, 22, 29, -17, -5, 21, 26, -1, 35, 2, 24, 19, 32, -18, 18, -13, -21, -11, -39, -17, -5, -23, -24, -21, -49, 1, -6, 37, 17, -10, -10, 16, 1, 40, 40, 21, 34, 21, -40, -12, 15, -27, -11, 6, 0, 45, 34, 15, -36, -22, -25, 11, -12, 12, 27, 33, -33, -29, 12, -29, 17, 46, 26, 7, 15, 7, -3, 48, 7, 13, -11, 21, 0, -31, -28, -21, -16, -32, 33, 13, 22, 1, -16, 1, 31, 41, -24, 31, -26, 36, 17, -28, 23, -25, -19, 33, 31, -25, -6, -14, 17, -5, 7, 14, -15, 20, 26, 3, 54, 22, -55, -42, -1, 44, -23, -66, -50, 11, -31, -67, -2, 3, 9, -27, 5, -26, 12, -7, 20, -29, 5, -5, -22, 3, 16, -36, -45, -14, 63, 45, 17, -9, 9, -6, -3, -8, -6, -15, 13, -27, 41, 2, -20, 13, -8, 14, -31, -2, -43, -47, 52, 33, 10, -32, 29, -6, -4, 28, -24, 14, -7, 22, -37, -3, -16, -30, -36, 41, 0, 51, 43, 21, 26, 46, 2, 56, -46, 3, -10, 7, 2, -45, 7, 4, 37, 41, 5, 62, -2, 13, 4, -36, -13, 26, -10, 25, 12, 60, 25, -5, -6, -36, 7, 1, 7, -18, -20, 13, -19, 17, -12, -5, 15, 16, 114, 26, 53, 23, 23, -19, 2, -30, -9, 47, 2, 39, 11, -1, -21, 21, 21, 42, -3, 0, -15, -35, -22, 45, 3, -27, -11, 15, 10, -8, 5, 39, 41, -5, 61, 13, -35, -47, 17, -5, 25, 11, -18, 21, -10, 41, -13, -4, 55, 48, 36, -34, -1, 6, -2, -55, -5, 7, 16, -23, -8, -5, -8, 25, -3, -39, 3, -12, 28, 3, -35, 6, -33, 32, -40, -24, -55, -46, -50, 28, 4, 10, -19, -39, -3, -22, -12, 17, -27, 34, 10, 19, -9, -50, -22, 7, -28, 5, 12, -21, 11, -41, 15, -19, -82, -18, 26, 43, -16, -6, -29, 6, 39, 23, 24, -78, 25, -26, 16, 27, 4, 0, -23, 11, 37, -4, -3, -19, 3, 35, -2, 13, 63, -14, 31, -33, 15, -49, 11, 14, -37, 6, 6, 15, 26, -23, 26, 39, 42, -21, 2, -27, 26, 19, 44, 4, 3, 9, -8, 50, -16, -37, -19, 34, 13, -22, 3, 35, -7, 23, 23, 35, -17, -12, -35, -29, 47, -4, 23, -26, -18, 5, 6, -9, -5, 13, 14, -10, 13, 25, -16, -15, 18, 19, -9, 28, 10, 20, -17, 1, -42, 3, -39, -4, -47, 1, -55, -24, -11, -18, -21, -18, -25, 23, 24, 22, 1, 44, 8, 30, 6, -23, -6, -6, 37, 33, 1, 22, 11, -30, -37, 13, -5, 3, -42, 22, -10, 21, -19, -6, 17, -8, 18, -16, 25, -31, 1, 13, -20, -44, -40, 28, 42, -16, 5, -5, -5, 51, -19, -26, 36, 47, 45, -17, 40, -21, 24, -39, 44, -31, -5, -23, 19, -39, 15, -11, 3, -28, -18, 20, 20, -4, 51, -6, -7, 60, 38, 4, 56, 2, -35, 43, -1, -41, 60, 17, 64, 41, -8, 41, -2, 14, 32, -19, 34, 36, 45, 32, 3, -3, 28, 36, 25, -21, 13, 14, 37, -67, 51, 53, 48, 0, 4, -27, -7, -21, 26, -10, -4, -41, -19, 24, 19, 7, 4, 6, 8, 23, -39, -36, 18, -19, -53, -31, 5, -4, -11, 13, 28, 25, 4, 24, 33, -24, -38, 20, -28, 42, -24, -44, 34, 18, 6, -22, -15, 8, 43, -7, 6, 19, 33, -12, 5, 36, 14, 16, 27, 29, 13, 12, 25, -5, 5, -36, -8, 27, -46, -53, -37, -21, -10, 39, 30, 28, 23, -30, -20, 33, -46, 29, 13, -42, -5, 38, 33, -7, -41, -32, 17, -20, 18, -18, -1, -9, -40, 8, -22, 21, 4, -28, -38, -15, 38, 27, 8, 1, 10, 39, -35, -19, -29, -48, 7, 24, 24, -4, -41, -41, 30, -40, -9, 32, 35, 41, -15, -3, 29, 36, 8, -8, 12, -1, 26, 6, 37, 12, -3, -26, -38, -34, 22, 25, 26, -30, -27, -7, 24, 41, -18, 4, 20, -29, 2, 27, -5, 9, 14, -15, 11, 61, 79, 17, -19, 29, -7, -31, 64, 56, 82, -2, -43, 2, 11, -8, 44, -29, 33, 18, -19, 11, 2, 30, 36, 38, 25, 1, 16, 21, 53, -2, -31, 3, 10, -14, 7, 25, -23, -28, 4, 40, -17, 30, -19, 22, -4, 2, 7, 15, -33, 43, -24, -27, -41, 12, -27, 34, -3, -12, -26, 13, 10, 17, 27, -6, 8, 26, 29, 39, -19, 32, -11, -46, -3, 19, -23, -9, -57, -12, -42, -7, 30, -24, -10, -39, -56, 32, -7, 7, -36, 9, -4, 11, 1, 4, 2, 6, -22, 22, -36, 23, -6, -40, -9, 14, 2, 4, 24, -6, 0, -12, 10, 9, -42, -11, -11, -10, 40, 5, -11, -18, 16, 18, -15, 16, 21, -38, 7, -55, 41, 41, -33, -13, 16, 30, -13, 5, -44, -10, 4, 14, -40, 23, 52, -41, 24, 31, 48, 34, 2, 13, -25, -7, -10, 24, 50, -23, 40, -20, 5, 17, -27, -26, 9, -26, 31, 7, -30, 30, -12, -4, -21, 22, -19, -4, -21, -35, -53, -21, 4, 38, -30, -21, 12, 38, -7, 30, 3, -34, -22, 32, 16, 28, -14, -37, -35, 5, -30, -41, -36, 7, -9, -28, 7, -25, -54, 82, 4, 19, -72, -42, 0, 30, -24, -34, 16, 31, -6, -9, -28, -58, 14, 17, 44, -78, -42, -54, 9, -11, -29, -4, -27, 4, 10, -23, -29, 34, 2, 18, -13, 37, 7, 8, -32, -49, -26, 25, -25, -7, -35, 1, -1, 28, -37, -23, -16, 12, 30, 30, 5, 24, 10, -11, -36, 6, 7, -14, -3, 27, -19, -26, 23, 41, -5, -36, -9, 13, -39, -15, 45, 0, 15, -9, 7, -7, 20, 36, -18, 15, 20, 12, 17, 22, -9, -3, 32, -19, 23, -12, 10, 5, -42, 37, 33, -18, 40, -33, -11, -17, -8, -41, -29, 4, -8, -5, -9, -39, -21, 41, -24, 7, 10, -7, -3, -32, -1, -1, 36, -7, -7, 3, -44, 12, 1, 27, -59, -21, -19, -29, 4, 13, -10, 37, 95, 14, -9, -4, 25, 9, 19, 36, -43, -4, 31, 34, 22, -12, 15, -25, 26, -30, 14, 3, 4, 2, -3, -23, 46, 12, -9, -44, -45, -35, 14, 26, 0, -9, -27, 6, -7, -32, -30, 2, -24, 18, -12, 19, 48, 6, 30, 14, 2, -9, -8, -7, -8, -13, 21, 29, -41, 12, 2, -1, 30, 46, 14, 26, 5, 37, 21, 71, 8, -25, 37, 33, 26, -17, -27, 17, -1, 19, 27, 8, -64, -11, -10, -3, -17, 0, 7, 43, 20, 18, -49, -8, 29, 58, 28, 40, 43, 54, 41, 4, 37, 36, -17, 15, -10, 17, -34, 10, -11, 29, -20, -13, 32, -35, 42, -13, 38, -2, -47, -14, -38, 0, -15, 22, 23, 31, 16, -27, -14, -41, -18, 7, 21, -15, 25, -11, 5, -36, -12, -30, -13, 32, -5, 34, 52, -23, -15, 13, 28, 8, 31, 26, -49, -28, -52, -40, -1, 29, 37, 32, -13, -22, 1, 15, 6, -19, -6, 37, 8, 13, -15, -48, 12, 26, -66, -64, 20, 44, 59, 29, 29, 19, 18, 55, -26, -24, -31, 12, -17, 23, -39, -13, 16, 36, 9, -13, -33, -14, 10, 61, 78, 24, -34, 24, -30, -24, -11, -9, 47, 42, 13, -26, 47, 17, 32, -7, -12, 45, 15, 32, -4, 34, 0, -21, -70, -52, 19, 16, 4, -14, -37, -34, 6, 35, 31, -21, 9, 38, 23, 41, -21, 6, 13, -3, 11, -35, -44, -4, -12, -14, -12, 2, 9, -8, -23, 8, 25, 26, -3, 10, -35, 18, 47, -12, -2, 26, 22, -25, -39, -5, 58, 54, -83, -58, -35, -39, -16, -37, -24, -25, -101, 45, -3, -50, -73, -39, -33, 7, 26, -21, 29, 49, 14, -2, 5, 79, 2, -23, -28, -22, -23, 8, -42, -29, -43, -9, -61, -18, 28, 48, 35, -51, 63, 1, 33, -45, -1, 27, 15, -9, 32, -5, 4, -14, -64, -49, -15, 19, 22, -43, -20, -3, 0, -5, -34, 1, -25, -35, 28, -22, -34, 6, -4, 15, 23, -17, -47, -52, 5, -12, 19, 37, 8, -28, 6, -43, -27, -1, 7, 20, -34, -23, 26, 29, 20, 27, -11, -22, 28, 0, 55, 18, -11, -22, 27, -36, 9, -36, -12, 15, 10, -21, -23, 32, 12, -40, -25, -22, -47, -14, 50, -33, 29, 21, -4, -39, -13, -25, 31, 11, -36, 13, 8, -28, -22, 16, 0, -35, 22, 63, -6, -27, -5, 27, -19, -14, 21, 30, 14, 13, -16, -35, -5, 1, -6, -51, 13, -13, 23, 0, -27, -1, 11, 13, 1, -22, 25, -1, -8, 20, 55, 34, -35, 24, -6, -8, 26, -29, 36, 15, 20, 36, 29, -46, -1, -8, -12, 0, -34, -12, -32, 2, -19, -20, 5, -3, 25, -28, 27, 18, 4, -55, 2, -25, 8, -5, 19, 28, -2, -27, 20, 21, 46, -23, -32, -9, -22, 9, -5, -8, -17, -9, 22, 47, -11, 32, -9, 22, 23, 21, 15, 37, -17, -22, 6, -46, -31, 15, 23, -2, -14, -8, -15, 55, 2, -6, -7, -20, -27, -13, 24, 4, 31, 26, 0, -15, 28, -23, -22, -36, 12, -31, -28, -4, -28, -2, 11, -38, 5, -2, 53, 7, 20, -12, 4, 39, 18, 9, 40, -20, -43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 24, -14, 35, -24, -29, -32, -16, -17, 21, -1, -20, -4, 50, 12, 14, -27, 30, 30, 21, -5, -10, -12, 37, 29, 25, 35, -5, -34, -13, 4, 26, -32, -18, -45, -16, -6, 15, 20, -25, 3, 7, 14, -29, 14, -19, 14, 0, 8, 54, 15, 13, 23, 4, 14, 16, 2, 26, 6, 40, -35, -14, 6, 36, -23, -1, 5, -15, -11, -7, 8, 36, -21, 37, 35, 2, 14, 55, 1, 15, 33, 38, -10, -43, -23, 20, 35, -5, 9, 12, 7, 50, 38, 30, 47, 10, 31, -19, 24, -14, 34, -30, -12, -34, 11, -45, -53, 4, 16, 1, -19, 4, 19, 52, -32, -16, 2, -5, 8, 26, -52, -8, -7, -18, 7, 11, 5, -23, -48, 17, 11, -41, -5, -48, -18, -32, 16, -8, 25, 43, -21, -14, -10, 8, -13, 30, 18, -41, 9, -49, 18, 45, 30, 11, -30, 8, -17, -36, -29, 6, -22,
 35, -1, -9, 33, 0, -55, 41, 21, 17, 26, 1, -31, 41, -4, 29, 27, 48, 48, -24, 3, 32, -37, 11, 28, 31, -31, -11, 36, -17, 14, 43, 19, 38, -22, -26, -21, 43, 39, -10, 27, 47, -11, 0, 4, -10, 7, -1, 22, -4, -23, 19, 3, -25, -22, 17, -21, 30, 15, 39, 29, 33, -23, 41, -21, 3, 69, 51, -12, -42, -12, 31, 58, -38, 12, 2, 25, 36, 29, 3, 4, -5, 24, 11, -8, 5, 27, 34, 51, 42, 10, 20, -8, 8, 15, 7, -6, -30, 23, -27, -18, 4, -4, 19, -3, 12, -18, 6, 38, 1, 2, 50, 8, -25, -24, 36, 31, -17, -60, 7, -7, 15, 36, 5, 11, -17, 19, 26, 15, 59, 17, -11, -26, -19, -7, 22, 13, -5, 24, -5, -1, 4, -13, 32, 27, 9, 22, 11, 19, -4, -23, 5, -5, 54, 9, -4, -3, -25, -1, 3, -1, -33, 3, -4, -35, -17, 7, 16, -13, 71, 4, -25, -12, 26, 52, 0, 43, 47, 46, 36, 4, 43, 31, -4, -10, -47, -40, -57, -12, -20, 4, 25, -4, -41, 15, -21, 0, -24, 17, 37, -30, 19, 3, -20, -35, 3, 40, 3, -21, -9, -2, 23, 14, 12, 10, 5, 28, -8, -45, -30, 20, 23, 9, -8, 23, 4, 38, -16, -3, -7, 21, 34, -31, 16, -11, 4, -11, 23, -19, 46, 22, 35, 26, 15, -32, -38, 10, -33, 36, 4, 37, -13, 29, 5, 34, -33, -37, -21, 18, -2, -46, 25, 5, -9, -24, 28, -15, -24, -35, 18, -10, -35, 22, -10, 21, 22, 26, 9, -36, -38, -62, 33, 36, 3, 10, -19, -45, 10, 20, 3, -11, -7, -33, -2, 29, -4, 10, 29, 6, 26, 4, 2, 45, -4, 26, -37, -24, -28, -16, -3, -53, -11, 31, -2, 18, -7, -24, -19, -25, -25, 13, -37, 1, 3, 31, -32, 17, -8, 4, -8, 5, 25, 23, 12, -2, 16, -36, -23, -36, -15, 35, 45, -4, -14, -23, -27, -19, -46, -27, 32, -33, -2, 13, 33, 30, -41, -8, -6, -71, -32, 118, 100, -18, -52, -58, -14, -10, 0, -40, -73, -17, 13, -22, -21, -7, 21, -33, -14, -16, 7, 41, 60, 25, -18, 7, -43, -37, -9, 33, 20, 20, 16, -19, 38, -19, -31, 7, -9, 38, 35, -40, 46, 46, 50, 4, -52, -37, -57, 3, 22, 11, -27, -4, -6, -7, -8, 37, 34, 32, 2, 18, 14, 11, 23, -36, -33, 22, 4, 21, 13, -55, -21, 35, -10, -33, 15, -6, -26, 14, -43, -3, 10, -12, -17, 7, -56, 11, 17, 0, 34, -40, 13, 19, -46, 13, -24, -9, 5, -15, 25, 8, 0, -6, 22, 35, 4, -2, 22, -1, 6, -27, -8, 26, 11, -20, -45, -16, -63, 20, 7, -34, 21, -38, -32, -6, -17, -26, -13, -4, -33, 11, 28, -27, -28, -44, -23, -48, 26, 10, -9, 2, -26, 30, -27, 0, -29, -9, 13, 21, -27, -50, -42, 42, 43, -13, -50, 35, -16, -6, -1, 4, 27, 24, 29, -29, -40, -5, -19, 6, -27, 31, 18, -41, -42, 11, 13, 17, 8, -20, 7, -34, -16, 11, -8, 8, -53, -31, 4, 41, 7, 27, 64, 26, -44, 11, 30, 46, 7, 21, 13, 9, 40, -18, -33, -10, -12, -3, -4, 6, -38, 27, 6, -10, 34, 27, -20, -22, -4, -41, -3, 29, 34, -47, -2, -34, 20, 44, 35, 3, 37, 13, -17, -17, -14, -37, -65, -9, 13, 25, 18, 11, 19, 1, -18, -44, 28, 22, -7, 32, 34, 16, -2, 46, 32, -5, -12, 39, 24, -15, 23, -5, 19, 21, 18, -24, -18, -8, 20, -30, -40, -29, 10, 29, -41, 40, 28, -37, 3, 43, -29, 12, 27, 38, 5, -5, -2, 32, 33, 26, 3, -10, -19, -14, -17, -11, -31, -6, -30, 7, -24, -6, 17, 14, 7, 27, 30, -17, 1, -15, -15, 12, 5, 33, 3, 5, -11, 8, -10, -3, 24, -33, -13, -18, -6, -2, -6, 26, -9, -61, -12, 7, 33, -21, -21, -15, 46, 28, -11, -13, -16, 6, -9, -9, -7, 2, -33, -3, 0, -19, 30, -2, 25, 13, -2, 28, 8, -14, -7, 9, 26, 11, -22, 24, -19, -6, -9, 5, 9, 14, 16, -29, -21, -14, -40, -20, -4, 18, 28, -1, -1, 21, 33, -16, -4, -6, 6, -13, -1, 17, 9, -48, -14, -38, -15, 0, 8, 11, 4, -42, -43, 10, 39, 90, 72, 45, -3, 7, -14, -35, -21, 16, 15, 11, -70, -42, 23, 31, 3, 3, -12, -43, -42, -39, -50, 31, -17, 14, 1, 4, -3, 39, 10, -5, -25, -1, 44, -1, 9, -26, -15, 5, -10, -10, -9, 12, -30, -2, -5, -23, 25, -1, 22, 22, 15, 19, 15, 15, 36, -17, 14, -5, -6, 50, 31, 3, -20, 15, 28, 5, 0, -25, -13, -16, -34, -2, -6, 21, -2, -12, 14, 12, 29, 11, 7, -43, -4, -37, 27, 10, -10, -26, 30, 33, 3, -8, -7, 46, -11, -16, -6, 14, 13, 38, 41, -17, 20, 42, -12, -18, 2, 9, -5, -11, -61, -68, -22, 32, -10, -7, 31, 28, -5, 17, -16, 56, 20, 33, -34, -33, -76, 29, 31, -10, -30, -47, -13, 14, 3, -17, 26, -9, 3, 38, -17, 11, 41, 45, 3, 9, 5, -4, 13, -21, 37, -56, 24, -26, 27, -45, -14, -38, -4, -4, -11, -22, -11, -1, -11, -13, 56, 9, -1, 24, -14, 46, 16, -1, 1, -8, -22, 24, 8, -57, -56, -28, -45, 1, 33, 34, 40, 26, -29, 1, 45, 40, -29, -6, -17, 11, -14, -70, -14, 100, -4, -65, 24, 24, -31, 7, 57, 15, -38, -24, 21, 56, -31, -33, -27, 61, 27, 7, -43, -67, 52, -17, -18, -6, 62, -2, 12, 21, -34, -27, -26, -16, 18, 15, 29, -21, 29, -1, -23, -4, -32, 16, 32, 4, -28, -40, 9, 15, -8, -37, 30, 12, 41, 12, 32, 30, -33, -12, 28, 36, -13, -16, -23, -19, 1, -33, 32, 3, 4, 18, -6, 16, 10, 14, -5, 16, -46, 38, 1, -37, -17, 7, 27, -4, 27, 28, -7, 12, 20, 42, 6, -11, -2, 9, -11, 21, -27, 5, 6, 5, 2, 19, 13, 16, 27, 24, 72, 9, 35, 26, 4, -68, 5, -21, 25, -36, -20, -30, 16, 36, 51, 57, 38, -44, 24, 55, -14, 17, 18, -31, 3, -15, 24, -37, -2, 21, -12, -31, -27, 37, 1, -66, 26, 9, -34, -17, 33, 1, -27, 6, 42, -6, -31, 50, 26, 53, 13, -27, 15, -17, 17, 5, 11, 23, 23, 43, 19, 33, -12, -19, 19, -22, 4, -16, -9, 3, -13, 19, 8, -18, -23, -10, 38, -6, -9, -9, -41, 54, -16, -23, 14, 19, 33, 40, -43, -2, 23, 18, 10, -58, -12, -33, 53, 23, 13, 36, 20, 20, 35, -7, -35, 41, 24, 48, 38, 37, 1, -12, -34, 25, -17, -32, 39, -24, -20, -35, -16, 24, -26, -3, -26, -12, -18, 3, 0, 12, -3, -44, -32, -2, -11, -18, -28, 9, -17, 18, -28, 18, -28, 20, 43, 36, 35, -15, 21, 40, -21, 6, -2, -6, 2, 10, 8, -9, 32, 4, -7, 28, 10, -3, 9, -26, -34, -17, 36, 11, -28, -18, 0, -35, 13, 37, -3, -44, 16, 32, -14, 15, 20, 31, -42, 18, 15, -20, -32, 13, 42, -30, -10, 13, 27, 32, -45, -28, 1, -3, 27, 10, -27, -15, -25, 25, 16, 31, -50, -38, -12, 11, -48, -23, 50, 31, -5, 27, -12, -4, -87, -21, 25, 16, 33, 39, -35, 12, 20, -30, 25, 20, 9, 20, -7, -49, -9, -9, -15, -42, 15, -17, 10, 11, 29, 27, -28, 6, 14, 30, 10, 20, -45, 15, 32, -16, -4, -38, 23, 31, 8, -12, -20, 16, -32, -16, 3, -22, 16, -39, -10, 18, -4, 13, 28, -16, 19, -20, -69, -47, -19, -20, -33, -15, 9, 24, 31, 33, 25, 11, -25, 10, 91, 15, 24, -30, 21, 21, 10, 7, 18, 29, -23, -12, -26, 23, -36, -3, 11, 18, -6, -5, 21, 4, -18, -33, -22, -20, 18, -15, 17, -26, 6, -14, -8, 15, 26, 7, 29, 25, -28, 8, 32, 44, -25, -4, -17, -2, -37, -46, 1, 12, 39, 19, 52, 10, -29, -37, -9, 7, 36, -11, -6, 23, -40, -13, -29, 2, -17, 13, -30, 7, 1, 12, 30, -11, 7, -27, 6, 11, 45, -21, -24, -3, 6, -25, -10, 14, -24, 30, 27, -3, 20, -9, 11, 8, 44, -13, 13, 3, -8, 33, 7, 24, 33, 8, 39, -22, 20, 56, 33, -10, -23, 29, 35, 4, -27, -13, -10, -48, -25, -16, -5, -27, 19, 33, 17, 18, 7, 6, 62, 32, 29, -21, 13, -48, -35, -3, 6, 36, 29, 7, -25, 6, 29, 20, -10, -34, -10, -26, -7, -19, -22, -9, -18, 31, 12, 34, 30, 6, 4, -15, 12, 32, 29, 14, -39, -32, -13, 17, -4, -11, -22, 42, 10, 14, -34, 11, 8, -3, 35, 5, 4, 23, 20, -32, 16, 18, 8, -11, -45, 78, 14, 53, 2, 35, -5, -32, 19, 15, 8, -14, -21, 11, 0, 34, 43, 32, -7, 8, -28, 8, -11, -48, -7, -21, -4, -20, 53, 33, 22, 8, 8, 20, 46, 14, -9, 29, 32, -18, 31, 16, 15, -11, -1, 3, 1, 23, 16, -34, 6, 3, 37, 5, 36, 13, 12, 16, -10, -42, -13, -35, -34, -47, -13, -6, -20, 2, 49, -11, 43, 25, 31, 17, -36, -23, 1, -13, -22, 26, -38, -37, -25, 54, -25, -24, -28, -27, -14, -27, -5, 11, -35, -15, -2, -9, 3, 33, -6, 42, -20, -4, 15, 1, 10, 9, -42, 23, 19, -23, -28, 26, -26, 23, -15, 3, 26, 31, 50, 62, 109, -20, -18, 2, 58, -22, -16, -24, -39, -9, -72, 29, -41, 8, -38, -32, 28, 0, -36, 16, 25, 18, -22, 33, 1, 45, 2, 23, -13, 37, 14, 17, -16, 25, 38, 11, 8, 19, 20, -36, 31, 27, 8, -2, -6, 19, -10, 9, 20, -10, -1, 14, -4, -35, -35, -36, -12, -25, -1, 9, 1, -26, -48, 29, -19, 11, 1, 15, 37, -19, -16, -11, -8, -5, 18, 38, 51, -1, -17, -20, -4, 78, 20, -29, -34, -1, 30, 30, 23, 20, -10, 27, 11, 0, 17, 34, 57, 55, -19, -47, 12, 66, 29, 6, -30, -7, 25, 10, -2, -1, 6, -28, -32, -10, -4, 16, 32, -45, -33, -15, 33, -1, -29, 24, -23, 40, -39, 1, 13, 31, -36, 21, -9, 30, 14, 8, -2, 15, 31, -30, -8, 1, -25, -18, 22, 33, 4, -11, 25, 8, 40, -39, 7, 20, 19, -11, 14, -5, 25, 25, 7, -5, -47, 18, -40, 29, -18, -1, 37, 18, -3, -43, 18, -20, 19, 36, -32, -27, -24, -5, 27, 24, 24, 41, 36, -9, 35, -31, -10, 3, 23, 37, 3, 34, -28, -5, -24, -16, -9, 23, -30, 30, -32, 27, 8, -10, 11, -12, -9, 45, 59, -11, 35, -34, 1, 53, -41, 41, 11, 18, -2, 27, 6, 27, 12, -2, 31, -10, -28, -5, -22, -18, -16, -6, 23, 16, 3, -30, -35, 43, -22, -45, -40, -23, -30, -5, -42, 5, 18, 3, -10, -38, -1, 1, -9, -32, 0, -10, 22, -16, 28, 41, 36, 27, 49, -21, -24, 7, -16, -15, 32, -21, 17, 53, 39, -18, -6, -7, -20, -19, -16, 0, 4, -10, 10, -11, -35, 67, -5, -39, -40, 35, 28, -9, -72, -10, 3, -49, 33, -3, -47, -54, -7, -14, -2, -13, -41, -47, -11, 17, 4, 17, 50, 27, -4, -21, 34, 31, 1, 13, 20, 16, 21, -25, 14, -16, 22, -22, 6, 18, 35, 26, 10, 45, 37, 31, 38, -5, -48, 15, -7, 18, 23, 18, 33, 24, -3, -30, 22, -32, 8, -40, 27, -12, 0, 30, -14, 49, -3, 41, 36, -2, -18, -29, -6, 27, 6, -22, -7, -27, 30, 22, 27, 22, 22, 28, 24, -13, 28, -1, -22, 51, -32, 11, 2, 15, -34, 24, -29, -21, -1, 0, 9, -28, -12, 33, 25, 16, -4, 13, -24, -5, 1, -5, 39, 3, 7, 1, -9, 61, 0, -27, 19, 20, -5, -26, 35, -10, 69, 17, 36, -6, -16, 44, -9, -19, 2, 13, 42, 30, -13, 32, -1, 6, 29, 25, -1, 39, 33, 28, 54, 15, -15, 46, -38, 10, 12, -21, -14, 13, 15, -21, 13, -9, 30, 21, -19, -27, 25, 20, 10, 20, -20, -34, -20, -48, 20, 18, 2, -9, 10, 12, 23, 33, 11, -8, 28, -21, 32, -4, -14, 2, 42, 3, -20, -36, -31, 16, -71, 0, -26, 34, -37, -29, -26, 9, 33, -3, -12, 27, -37, -14, -41, 45, 33, 15, 22, -27, -33, -25, -34, 10, -25, -5, 18, -21, -53, -22, 22, -31, -11, 32, -16, 8, -7, -24, 39, 13, -13, -19, 22, -23, -13, -2, 54, 31, 25, -4, -8, 55, 25, 20, -15, -1, 0, -7, 0, -29, -22, 18, -8, -7, -26, -3, -11, 5, 7, -28, 11, 26, -15, -31, -38, -6, 37, -38, -32, -38, 16, 6, 35, 9, -5, 2, -14, -52, -9, 4, -4, 19, -18, 9, -17, 7, 34, -29, 6, 17, -10, 13, -37, 0, 38, 0, 3, 20, -25, 15, 45, -28, -51, 16, 18, -5, -9, -72, -2, 12, 20, 2, 8, 24, 19, 17, 25, -10, -7, 29, 4, 30, 56, 15, 4, 2, -56, -67, -8, -6, -13, -22, -34, -5, -8, 41, -32, -70, 10, -35, -1, 0, 6, 7, -12, 9, -30, 10, 2, 35, -3, 4, -62, 15, -14, 40, -43, -68, 11, 37, 28, 13, -43, 21, -3, -12, 7, -34, -11, -12, -1, -24, 28, 10, 20, 35, -34, -57, -25, 5, -6, 52, -45, -13, 27, 3, -37, 15, -29, -15, 4, 12, 16, 19, 27, 20, 33, 4, 28, 33, -40, -115, -81, 20, 16, -18, -27, -57, 7, 14, 1, 2, -88, -5, -31, -39, -26, -41, 3, 49, 10, 11, 40, 21, 35, 12, -18, -78, 15, 19, 51, 23, -73, 15, -12, 6, -19, -43, 13, -28, 21, -19, -26, 12, -2, -15, 38, 25, -8, -17, 23, -46, -74, -13, -27, 50, -12, -72, -17, 39, 26, 36, -23, 36, 7, 24, 5, 16, -14, -14, -1, -6, 2, 10, -18, -31, -28, -15, 21, 35, -21, 38, 44, 9, 40, 28, -44, 38, -21, 32, -30, 37, 36, 14, -22, -31, 16, -11, 1, 60, 50, 62, 78, 30, 11, 10, 32, 41, 5, -33, 37, 54, -42, 41, 27, 0, 3, 16, -11, 27, 40, 22, -40, 1, -13, 3, -21, 56, 15, -24, 13, 64, 16, 35, 58, 38, 32, 19, 33, 30, 26, -32, 25, 18, -5, 28, -13, 9, 0, 78, 18, 4, 16, 9, 15, -2, -19, -29, -34, 21, -32, -29, -4, -16, -20, -27, 22, 29, 1, -4, -20, 26, -29, 35, -27, -39, -23, -7, 24, -7, -19, 8, -4, 25, -23, 1, -60, 24, -39, -36, 9, -15, 6, -36, -35, -38, 5, 3, 49, -18, -52, 0, -58, 1, -49, -76, -20, -41, -22, -29, -31, -18, -41, -23, -22, -19, -7, 42, -48, -40, -10, -12, -17, 3, 2, 25, 29, 24, 22, -6, 40, 48, -17, 1, -5, 8, -41, -19, 41, -4, -19, 22, 14, 19, 21, 16, -28, -50, 44, -2, 32, -12, -1, 13, 6, -22, -9, -34, 26, 12, -13, 8, 18, 25, 17, -46, 19, 26, -19, -31, 41, -31, -39, -17, 10, -14, -8, 21, 13, 8, 27, -25, 0, -7, -2, 20, -38, -17, -43, -13, -22, -15, -43, 38, 25, 20, 21, -13, -34, 40, 27, -22, -34, -38, 18, 4, -16, 13, 18, 24, 27, 19, 38, -34, -12, 41, 27, -23, -25, 4, 19, -8, -1, -18, 18, -2, -26, -6, 6, 26, 33, -22, 24, -20, -44, -7, -43, 14, -5, -28, -14, 16, 31, -11, 19, 10, 33, -20, 14, 27, -14, 39, -22, -4, -36, 0, 26, 31, -29, 18, -2, 8, -5, 11, -22, -18, -29, -31, -20, 0, 13, 4, -30, -10, 24, 9, 0, 23, 29, -49, -17, 37, -12, -29, -7, 28, -16, 7, 39, 13, -20, 37, 1, 24, 99, 52, 3, 1, -8, 31, -9, 9, -34, -1, -18, 5, 32, 44, 43, 50, 27, -31, -11, -19, -7, 23, -34, -51, 14, -5, -57, 6, -21, -10, -19, 45, 38, 38, 22, 10, 14, -36, -12, 7, -46, -21, 23, -3, 10, -40, -44, 24, 18, 8, -11, 19, 14, -36, 14, -9, 44, 26, -28, -24, 19, -12, -14, -21, -28, -5, -22, -2, 9, -20, -30, 1, -22, -36, 35, -37, -29, 6, -33, 12, -2, -16, 17, -20, -14, -8, -22, -26, 5, -36, -1, 0, -8, 20, 3, -19, 2, -4, 11, -11, 2, 26, -11, -2, -27, -67, -2, -44, 17, 5, -39, 14, -25, 59, 16, 14, 29, 1, -44, 30, 4, -2, 0, 27, 10, -28, -31, -38, 34, -18, -11, -10, -34, -6, -3, -20, -32, -18, -11, -20, -20, -32, 33, 14, 10, -4, -5, -26, -19, -16, -21, 6, -9, 32, -26, -2, -4, 16, -7, 8, 16, 30, 21, 4, 2, 24, 25, -5, -18, 25, 6, 25, -15, 15, 6, -7, -19, -17, -1, 8, 7, 39, 36, 10, 24, -8, 31, 12, 24, 14, 24, 39, -11, -18, 72, 19, 26, 43, 0, 20, 6, 9, 32, -10, -19, 46, 20, 26, -20, 38, 17, -5, -19, -25, 28, 32, 32, 43, 43, 1, 25, 39, 0, 18, 17, 3, 3, -23, -12, -7, -15, 27, 13, -1, 5, -12, -19, -13, -47, 28, -26, 30, 46, 36, -31, 0, 20, -24, -22, -18, 28, -4, -15, 7, -1, -39, -2, -6, 1, -6, -16, 37, 8, -30, 6, 15, 16, 9, 14, -17, 6, 30, 1, -13, 6, 7, -1, -2, 8, 28, -15, -25,
  1, 19, -15, -2, 30, 4, 17, -17, -18, -24, -27, -9, 40, 18, 32, 17, 1, 43, -8, 22, -3, -7, -33, 10, 23, 33, 2, -36, 20, 31, 33, 28, 20, 23, -42, -15, -10, -37, -40, 51, -4, -1, -7, -8, -19, 20, 23, 23, -19, -9, -19, -41, -40, 31, -13, -46, -43, -12, -2, 13, 2, -15, 28, 56, 38, 18, 1, 28, 40, 26, -12, 31, -2, 9, 10, 28, 6, -34, 23, -17, 7, 51, -25, -25, 9, -3, -44, -3, -21, -14, -51, -54, 34, 17, 26, -9, 57, -29, 5, 23, 16, 7, -13, -22, -37, 5, 20, 39, 24, -13, -75, -34, -15, -64, -54, -34, -17, 1, 13, 48, 24, 63, 3, 14, 27, 29, -34, -15, -1, -1, 55, 0, -31, 40, 0, -14, -57, -25, -42, 7, -42, 16, -10, -20, -11, -25, 35, -19, -5, -3, 36, 27, 13, -29, 24, 33, 19, 27, 31, 16, -10, 9, 13, 21, 37, -37, 17, 31, -10, 24, -11, 17, -18, 39, 5, 30, 22, -23, 5, -13, -8, 43, -10, -36, 1, -40, -34, -40, -18, 26, -11, -12, -13, 14, -16, 4, 38, -20, 10, 7, -4, 9, -6, -19, -31, -7, -12, -41, -29, 29, -5, -32, -27, 17, 50, -22, 40, 13, 38, -23, -33, -10, -35, 10, 3, 70, 78, -25, 12, 35, -10, 29, -4, -23, -7, 22, 12, -11, 33, 69, -28, -25, 14, -28, 6, -10, 25, -34, 5, -36, -21, 26, -31, -29, -27, 15, 2, -39, 22, 37, 26, 60, 49, 52, 30, 4, -15, 12, 1, -17, -1, -27, 24, 16, 21, 37, 15, -5, 29, 40, 15, 22, 2, -35, 8, -3, -16, -16, -43, 31, -27, 12, -12, -18, 13, 29, 24, -9, 40, -50, -35, 23, 29, -6, 16, -4, -6, 67, 67, -5, -23, -55, 33, 0, -29, -3, -8, -27, -41, -11, 57, 66, 16, 75, 30, -8, 14, 13, 7, -42, 10, -27, 36, 21, 29, -16, -6, 4, 11, 33, -9, 34, -17, -3, 9, 9, 7, -26, -17, 36, -10, -32, 34, 26, 7, -18, 38, -9, -21, -35, -5, 28, 46, 55, -17, 24, 17, -10, 21, -39, -44, 33, 14, -1, 25, -8, 38, 39, -32, -21, -29, 41, -27, 12, 34, -20, -28, -33, -16, 54, -41, 4, 22, 16, 13, 39, 13, 19, -23, 37, -14, -28, 0, -16, 6, -8, 50, 0, 25, -12, 40, 12, 10, -28, -14, 33, -19, 26, -17, -7, -26, 13, 7, -30, -71, -12, -25, -46, 15, 0, 8, -10, -45, -36, 14, -30, -7, 35, 4, -22, -8, 39, 15, -32, -17, 25, -38, -21, 28, -19, 33, -48, 20, 20, 27, -16, 10, -49, 23, 11, 39, 14, -29, -14, -18, 29, 28, 18, -18, -24, 7, 18, -4, -47, -11, -5, -11, 11, 18, 15, 8, -6, 1, -42, 27, -16, -12, 34, -4, -6, -23, 38, -9, 15, -18, 26, -22, -28, 27, 42, 7, -15, 59, 13, -2, 24, 54, -13, 18, -39, 17, -24, 14, 55, -2, 32, -8, 4, -25, -20, -40, 2, -7, -3, -7, -16, -18, 34, 31, 18, -3, 30, 16, -22, 28, 36, -2, -10, -1, -36, -17, 9, 34, -21, -32, 34, 24, 21, 26, -36, 49, -5, -13, -1, -17, 28, 15, 11, 41, 57, 11, 7, 40, 30, -3, -19, -3, -21, -21, 18, 22, -25, 1, 25, 31, 2, -25, -5, 3, -29, 26, 34, -30, -48, 35, 40, 23, -21, 26, -11, -26, 9, 36, -41, -38, -25, -15, 4, 15, 12, 9, 47, -17, -30, 1, 57, -11, -2, 35, 13, 19, -10, 5, -16, -14, -2, -36, -12, -27, 19, -35, -53, 1, 13, 14, 27, 2, 1, 38, 18, -10, 40, 13, 57, 17, 8, -2, -47, 18, 6, -5, 15, 10, 15, 39, -2, -67, 25, 20, -28, 31, 41, -21, 15, 31, 6, -1, 23, -5, 41, 30, 24, -20, 18, 15, -39, 4, -24, 10, 19, -1, 40, -28, -26, -4, 62, 3, 38, -27, 2, -25, 23, 2, 2, 44, 34, -13, -46, 4, -18, -13, -13, 33, 18, -1, -35, -20, -5, -14, -14, 24, 15, -54, 2, 0, 30, -26, -46, 4, 40, -2, -49, -28, -51, -63, -26, -33, 30, 25, 27, 45, -30, -25, -30, -12, 16, 12, 45, -28, -14, -32, -27, -35, -64, -2, 21, 6, -49, -36, 16, 34, -31, 23, -44, -9, -53, -30, -24, -13, 13, -8, 49, 18, -43, 30, 35, 32, -30, -16, 17, 55, 18, -52, -21, -15, 16, -43, 25, -17, -31, -15, 4, 43, 6, 34, -2, -20, 38, -15, -12, 32, 0, 15, -10, 20, 30, 6, -7, 23, 2, 5, 20, -12, -35, -5, -20, 3, 27, 9, 15, -24, -22, -34, -22, 15, 20, 17, 38, 46, 2, -37, 47, 19, 35, 26, 6, 39, 47, 3, 3, -35, 5, -11, -29, 64, 59, 63, -31, -29, 33, 62, 56, -26, -8, 19, 46, 21, -27, 8, 9, -8, -16, 14, 18, 3, -18, 31, 34, 10, -16, 30, -16, 12, 18, 3, 39, 11, 31, 49, -22, 2, 46, 4, 18, 10, -1, -25, 36, -18, -48, 16, -47, 22, -27, 7, 43, 33, -5, 43, 3, -7, -33, -5, 37, 30, -40, -1, -39, -5, -10, 23, -10, 5, 47, 27, 35, -3, 9, 7, -1, -19, -31, -36, -41, 10, 20, -12, 7, -6, -8, -21, -11, -22, -50, 11, 7, -31, -57, -21, 24, 15, 42, 35, 8, -43, -40, -39, 18, -26, 0, -14, -68, -10, -20, 19, -55, -12, -24, -41, 0, 7, 54, 7, -30, -5, -7, 35, -16, -38, 23, -13, -19, 5, 27, 10, 7, -12, -4, 26, -22, 33, 29, 29, -29, -4, 29, 27, 8, -5, -42, -25, -8, 5, 4, 29, 1, -38, 3, 31, -3, -8, 28, -7, -25, 21, 8, 7, 35, 33, 13, 17, 24, 17, -14, -19, 22, -16, -10, 25, 35, -8, 41, 20, 11, 6, -46, 11, -18, 9, 45, -11, 36, 33, -7, 22, 14, 7, 4, 33, 13, 5, 22, -34, 21, 55, 65, 110, -34, -7, -28, 27, 55, 18, 21, 5, -5, -68, 29, -10, 3, -44, 45, -10, 12, -21, -12, 3, -26, -30, -4, -7, -36, -1, -39, 20, -9, 42, 14, -46, -6, 11, 36, 16, 3, 32, -42, -70, 40, 39, 28, 7, -8, 10, 41, 42, 37, 7, 34, -19, 24, 9, -45, 30, -29, 51, 5, -6, -18, -23, 8, -5, -30, -15, 12, -31, 9, -1, -11, 52, 26, -9, -18, 6, 19, 17, -27, -13, 9, 56, 33, 23, -1, 76, -23, 25, 32, 8, -18, -5, 24, 35, 1, -10, 56, 50, -47, -6, 49, 19, 6, -52, -6, 55, 24, 41, -6, 64, 30, 21, 26, 41, -5, 19, -10, -12, -22, -42, -17, 28, 15, -46, -32, -22, -47, 1, -25, 19, 0, -25, 15, 3, 4, -33, 24, -21, 8, -30, 34, 34, -51, 15, 14, 24, 5, 8, 31, -9, 5, 32, 32, 32, 11, -8, -2, 44, 24, 6, 0, -41, 36, -42, 3, 30, 9, 15, 25, 11, -21, 20, 9, -48, -83, 38, 5, 43, 25, -47, -5, 1, 17, 1, 5, -40, 32, 1, 44, -12, -49, -35, -16, -12, -38, 8, 15, -60, -48, -59, -15, -21, -36, -13, -2, -11, 9, -5, 39, -17, 29, -18, 10, -16, -41, -23, -11, -7, 35, 10, 8, 47, -1, -38, -44, 56, 1, 15, -44, -43, -18, -37, -3, 56, 17, -23, 13, 8, 13, 22, -23, 21, 3, -28, -32, 31, 13, -25, -66, -57, 29, -14, 45, -19, -39, 30, -31, 8, 37, -17, -42, -20, 42, 16, 10, -22, 26, 19, -37, 13, -20, -8, 25, 14, -38, 61, 26, -3, 58, -12, -22, 2, -42, 9, 28, -9, 21, -6, 1, 26, -32, -40, -50, 10, 0, 24, 39, -20, -64, -76, 23, 28, 28, -4, -12, 10, -29, -38, 23, -67, 22, -37, -13, -16, 41, 6, -31, 4, 0, 32, -3, -12, 27, -57, -58, 23, -16, 36, 4, -25, -9, -33, 36, 51, 19, -21, 18, -12, -2, -18, -5, 22, -27, -38, -50, -4, 42, -30, -64, -24, 30, -30, 29, 8, -27, 36, -31, -10, 37, -10, -47, 22, 11, 31, -13, -49, -46, 46, -31, -25, 25, 29, -27, 4, -34, 23, -21, 18, 27, -5, -37, 11, -7, 25, -16, 15, 24, -2, -39, 13, 22, -26, 23, 28, 45, -18, 40, 33, 57, 51, -6, 9, -5, -8, -67, 22, -8, -9, 17, -31, 33, 15, 22, -11, 36, -10, 18, -51, 11, 27, -1, -16, -24, 39, 31, 21, 24, -18, 32, -21, 3, 30, 38, -22, 12, -23, -10, 35, -9, -48, 1, -33, -4, 2, -11, 49, 11, 14, 2, 44, 8, -5, 27, -30, 8, -17, -34, 34, -2, -16, -10, 4, -4, 2, 9, 12, -20, 15, 23, 29, -36, 23, -6, -31, -50, 44, 19, 9, 22, -25, 50, -41, 34, -23, 19, 52, -41, -15, 28, 56, 41, 49, 0, 13, 37, -9, 35, 32, -27, 32, 38, 21, -10, -46, -54, 2, 6, -7, -13, 16, -5, -43, 40, 12, -9, -10, 24, 27, 52, 34, -12, -33, 8, -19, -4, -4, -4, -30, 28, -21, -5, -4, -2, -20, -15, 1, -4, 20, -2, -6, 2, -15, -28, 41, 14, 2, 22, -7, -12, -1, -5, -42, 25, 14, 15, 16, -10, 10, -17, 27, -1, -16, -3, -41, -1, 36, -11, 35, -28, -6, 5, -17, -27, 27, 35, -4, 10, 32, 14, -1, -21, 16, -30, -30, -16, -12, 40, -8, 0, 10, 10, 9, 21, -11, 17, -3, -4, 31, -21, -61, 5, -9, 8, -14, -12, -18, -14, 39, 31, 19, -11, 46, -9, -5, 31, 47, 47, 15, -32, -55, 3, 46, 25, 23, 22, 4, -23, 15, -30, 21, 19, 39, -20, -5, -18, -3, -2, -2, -32, -2, 35, 13, 3, 8, -21, -29, -24, -34, -21, 8, 30, -3, 22, 26, 32, -2, 2, 49, 13, 21, -8, -3, 6, 43, 6, -15, 32, -19, 15, 11, -37, -15, -20, 22, 14, -55, -44, -12, 1, 48, -56, 19, 8, 40, -12, -30, -48, 2, -22, 34, -14, 26, 82, 46, 35, -50, -22, 4, 33, 42, -71, -5, 32, 57, 13, -46, -4, -6, -13, -20, 2, -19, -14, -19, -45, 23, 15, 36, 1, 9, 5, -32, 43, 25, -26, 10, -21, 32, 10, 31, -18, 31, -22, 7, 7, -15, -7, -10, -37, 19, -4, -13, 13, 30, -27, 8, 27, 4, 38, 13, 38, -27, -9, -34, -4, 29, 31, 17, 14, 38, 19, -10, 5, -24, 36, 35, -3, 7, 23, 0, -22, -19, 20, 16, -26, -53, -20, -4, 5, 7, -45, 29, 7, -1, -23, 19, -22, 32, -19, 6, 40, -5, -16, -29, 36, -8, 23, -35, 41, 50, 16, -42, 5, 87, -1, -11, -53, -38, 35, -53, 19, 19, 22, -59, -15, -25, -28, -14, 34, 7, 13, 22, 19, 9, 9, -24, -8, -8, 21, -4, 1, 40, 44, 0, -39, -21, 8, 39, -30, -45, -4, 6, 14, 10, -53, -31, 18, 24, 10, 35, 9, -30, 1, 6, -27, -29, -61, -33, -5, -46, 18, 3, -29, -14, -15, 12, -23, -26, -15, 10, 50, 61, 10, 48, -9, 26, 33, -7, -46, 3, 45, 26, -32, -10, -15, -7, 4, -19, -27, -4, 13, 41, 16, 25, 4, 30, 48, 26, 8, -37, 88, 39, 9, -20, -64, -10, 46, 1, -34, 1, -1, 9, -29, -11, 0, -29, 41, -3, 32, 29, 2, 41, -36, 35, 16, -48, -31, 16, 22, -24, -29, 3, 6, 32, -35, 49, 49, 6, 46, 6, -24, 12, 7, -3, 24, -13, -20, 11, 35, -24, -4, -43, -34, 55, 14, -54, -19, -18, 34, 1, 5, -19, -8, -34, -20, 4, -37, 31, 41, -20, -20, -17, -14, -15, 0, -10, 25, 23, -11, 6, -45, -40, 17, 12, -14, -40, -52, -35, -9, -2, 32, 33, -21, 57, -18, 1, 26, 1, -2, -12, -31, -39, 43, -35, 1, -45, 28, -24, -6, 18, -16, -33, -1, 40, -5, -16, -38, -7, 31, 22, 31, -17, 28, 28, 3, 30, -21, 3, -38, -21, -49, -19, 21, -59, 13, -38, -21, -9, -24, 6, -27, -60, 10, 22, 3, 32, -14, -16, -26, -19, 31, 2, -33, -15, 11, 9, 16, -3, 1, -7, -29, -51, 38, -1, 60, 44, -15, 21, 24, 22, 38, 51, 46, 20, -24, -7, -16, 9, -57, -70, -29, -37, 39, 6, 30, 31, 71, 4, 11, 4, 49, 70, 44, 43, 20, 38, 3, 22, 13, -19, -3, -21, 16, 51, 7, 2, 30, -14, 20, -50, -14, -1, 13, 19, 33, 38, 0, 33, 28, 28, -27, 16, 37, 11, -7, -8, 9, 9, -27, -45, -24, -26, -16, -30, 20, -24, 0, 8, 32, 5, -31, -8, 53, 24, 3, 15, -21, 30, 21, 5, -7, -1, -18, -46, -52, -50, -41, -12, -21, -35, -20, -6, 22, 43, 5, 13, -40, -9, 23, -6, 8, -26, -6, -32, -32, -4, 5, -3, -9, -26, -4, 0, -7, -15, -28, 12, 6, -29, 38, 5, 35, 29, 3, -15, 37, 6, 5, 31, 30, -2, 16, -16, -32, 71, -21, 24, -10, -48, 40, 42, 2, 15, -7, -9, -13, 23, -4, 34, 7, 43, 1, 22, 8, 27, 17, 14, -23, -3, 60, 30, -30, 41, 27, 32, 19, 5, -22, 43, 30, 73, 38, 31, 20, -34, 1, 28, 13, 40, 32, -34, 20, 19, 2, -20, 9, 17, 14, -8, -7, -48, 27, 19, -25, 12, -38, -8, 19, -8, 38, 16, 33, -10, 1, -22, 2, 38, 39, -23, 4, -20, 81, -29, -51, -59, -37, 10, -22, -13, 12, -6, 14, 31, -37, 17, 7, 42, 1, 1, 11, -39, 61, 26, 26, -41, -45, 5, 43, 51, -21, -29, -1, 0, 17, 13, 16, -9, 36, 2, 25, 26, -26, -9, -7, -6, 9, -26, 20, 49, -1, 39, -8, 15, -27, 33, 14, -16, -21, -4, 22, 42, 18, -31, 27, 1, 4, -38, 33, 42, 51, -18, 17, -7, -28, -6, 24, -34, -34, -26, -11, -33, -36, 3, -33, -11, -13, -15, 23, -32, 19, 39, -27, 2, -19, 3, -47, -22, 17, -40, -36, 29, 11, -8, 34, 13, 3, 37, 2, 26, -20, 37, 12, 1, -31, 19, -23, -43, 45, 95, 62, 18, -7, -23, 68, 0, -58, 6, 11, 29, 19, 21, 28, 18, 38, 40, -27, -1, 19, -10, 13, -19, -18, -40, 17, 5, -5, -25, -23, 40, -27, -19, 6, -15, 23, -11, 30, -9, -36, 45, 12, -15, 14, -11, -18, 8, -24, 11, 24, 15, -3, -61, -23, 12, -22, 4, -75, 8, 23, -29, -28, 40, 24, 3, 16, 42, 56, 33, -15, -31, -29, -3, -8, 17, -49, -20, -18, -1, -41, -37, -15, -25, 26, -22, 53, 30, 27, -17, -18, -12, -23, -8, -8, 12, 20, -13, -36, 2, 48, -1, 5, 44, 8, -13, 1, -50, 4, -4, -20, 32, -13, 30, 47, -17, -23, 20, 71, 16, -9, 18, 25, 8, -4, -23, 36, -42, 6, -20, 12, -19, -31, 18, 35, 47, 44, -14, -9, 4, 12, -39, 26, 23, -26, -44, 30, -37, -9, -24, 25, -10, -19, -31, -23, 10, 0, -62, -28, -17, -6, 7, -18, 31, 28, -48, -5, 43, 29, -13, -14, 12, 27, -4, -4, 43, -15, 21, 23, -35, 1, 8, 35, 0, -7, -38, 37, 1, 7, 19, -33, 7, -31, 8, -16, 10, -24, 8, 10, -28, 5, -17, -16, 23, -12, -51, -49, 49, -5, -41, -47, -35, 18, -65, 0, -27, -11, -18, 3, 17, 22, 15, 6, -12, 5, 13, 17, -17, -5, -40, -12, 3, -29, 32, -11, -29, 27, 17, 3, -32, 0, 43, -4, -55, -28, -11, 3, -43, -15, 34, 38, -3, -1, 34, -12, -16, 4, 48, 30, -3, 1, -37, 19, -43, -64, -11, 9, -25, -7, -28, -7, 6, 30, -20, -1, 16, 3, 41, 10, 18, 34, 21, 23, 14, 79, 42, -45, -19, -39, 34, -48, 39, 14, 62, 34, 15, -12, 20, -8, 29, 30, -10, -5, -8, 8, 52, 70, 36, 13, 26, 47, -25, -9, 7, -32, -30, 9, 25, 1, -27, -3, -5, -16, 14, 18, -7, 13, 0, 27, -9, -41, -35, 26, -16, 5, 24, 20, -2, -15, 9, -28, 30, -21, -42, 23, 31, 4, 13, 4, -19, 15, -13, -10, -2, 6, -5, 18, 10, 39, -47, -18, 0, -14, -42, -2, 7, 4, -45, -37, 26, -31, 32, 28, 27, 26, -18, 23, 12, -4, 15, -20, 35, -17, -28, -44, 1, 8, -3, 41, 31, 29, 41, -19, 24, 18, 35, 13, -13, 29, -12, -28, -19, -30, -54, -13, -62, -47, 14, 32, -26, -29, 26, -60, 12, -20, 4, 5, 15, -45, 32, -2, -35, -2, 17, -19, 10, 19, -9, -75, 5, -21, -3, -21, -40, 7, 9, 36, 25, 0, -15, -15, 10, 5, 8, 21, 2, -46, -25, -34, 30, -30, 13, 9, 49, -30, -49, 25, 5, 42, 33, 10, -1, 18, 35, -26, 15, 16, 32, 41, 13, 13, 36, 37, -7, 8, -9, 19, 31, -34, 48, -2, -26, 17, 21, 27, 33, 37, 19, -19, -18, 17, 34, -13, -26, -11, 16, 73, 21, 1, -28, 22, 13, 0, 21, 2, 27, 36, 30, -12, -9, 21, 59, 24, 19, 12, -37, 54, -16, 28, 26, 36, -1, 14, -27, 10, -27, 36, 2, -3, 29, -18, -2, -45, -44, -4, -23, 1, 7, 4, 14, 3, 21, -10, -30, -5, -6, -45, -12, -2, 18, -34, -19, -4, -20, 12, -41, 5, 25, 32, -8, 3, 18, -6, 25, -30, -22, 49, 26, -7, 39, 2, -9, 40, -44, -6, 35, 43, 21, 51, 20, -35, 14, -28, -16, 14, 14, 16, -39, 22, -14, -37, 2, -20, -37, 9, 20, 33, -10, 57, 18, -5, -38, -21, -17, -15, -19, -40, -30, -44, 9, 24, -18, 9, -64, -48, 34, 32, 5, 17, -3, 16, -28, -35, 1, 27, 27, -19, 14, 4, 32, -6, 11, -2, 33, 35, -11, 3, -15, -63, -2, -1, 25, -20, -30, -35, -7, -29, 77, 5, -29, 27, 29,
   9, -29, 28, -4, -15, 37, 6, 6, 31, 9, -4, 17, -4, -19, 52, -13, 28, -52, -46, -42, -17, 26, -28, 56, -8, 31, 6, 28, 12, -22, -5, -11, -14, 12, 9, -22, 4, -33, -80, 10, 28, 28, 43, 21, 50, 62, 73, -41, -20, -38, -52, -31, -2, 46, 48, -7, -8, 3, -20, -39, 15, 57, -18, -21, 22, -24, -92, -26, -18, -12, -2, -10, 8, 38, 40, 49, -26, 19, 0, 39, 29, -3, 6, -20, -12, 22, -12, 2, 5, -42, -19, -22, -38, -14, -7, 14, -7, 24, 36, 38, -6, 11, -6, -43, 8, 26, 29, 1, -25, 53, 15, 37, -21, -39, 7, -25, 36, -18, -21, -11, 19, -7, 24, 14, -24, 4, 28, 35, 18, 40, -14, -11, -18, 22, 42, -16, -12, -11, 30, -11, 2, 14, -17, -27, 19, 21, 2, -6, 12, -71, -54, -23, 13, 3, 3, -7, -64, -34, 30, -28, -27, -13, -27, 32, -47, -5, 33, -30, -44, -7, 43, 35, -13, 14, 1, 26, -16, 22, -18, 18, -19, -16, -34, -13, -21, -32, 9, 7, 38, 6, 9, 8, -24, 13, 10, 35, 42, -16, 2, -40, -43, -53, 30, -14, -29, 15, 3, -20, 21, -35, -18, 29, -25, 18, 3, -6, 27, -23, -45, -18, 7, 18, 15, 57, -1, -25, 12, 20, 55, 27, -30, -16, -12, -9, 25, 28, -8, -11, 10, -28, 23, -1, 58, 6, 5, 0, 19, 11, 32, 7, -42, -6, 9, 42, 25, -21, -32, 23, 28, 0, -23, 13, -3, 60, 41, 21, -27, 2, 24, -1, -2, -38, 7, 13, 3, -1, 5, -24, 25, 0, -17, 24, -12, 44, 7, -20, 10, -27, 52, 11, -25, 31, -31, -2, -22, 6, 41, 6, -8, -11, -36, 11, 30, 15, 31, -17, -34, -10, -22, -1, -25, 13, 19, 32, -1, -18, 0, -34, -19, -1, 12, -7, 18, 26, -9, 4, 14, 31, 11, -24, -13, -2, 37, 19, -34, -11, -9, 34, 6, -23, -29, 9, 5, -11, -1, -16, 0, 12, -29, -20, -22, 23, 24, -18, 6, -6, -11, 16, -17, 18, 2, -2, 18, -13, -28, -3, 23, 7, -1, 5, 14, 2, 20, 1, -6, -2, 2, 21, 8, -13, 0, -5, 23, -35, -33, 5, -24, 25, 0, -15, -19, 19, -3, -18, -32, 13, 41, 12, -29, -36, -27, 5, 16, -3, -21, -6, -22, 22, -15, 13, -6, -6, 17, 2, -34, 5, 11, 11, 12, 6, 16, 11, 21, 17, -7, 14, 7, 37, 31, 0, -9, 0, 10, 17, 19, -10, 1, 22, 27, 4, -5, 8, -18, -23, 0, 19, 19, -34, 2, 19, 2, 25, -3, -8, 22, -12, -11, 19, 13, 23, 19, 41, 10, -5, -18, -10, -20, 7, 20, 1, -10, 18, 16, 19, -25, 4, -8, 17, 18, -5, -11, 3, 20, -3, -18, -4, 5, 25, -10, -15, -19, -9, 0, -7, -13, 19, 36, 19, -15, -2, -14, 4, 25, 3, -9, 11, -11, 24, -1, -6, 3, -13, 22, 2, -21, 0, -1, 6, -23, -3, 2, 3, 36, 19, 22, -21, 23, -3, -29, 26, 5, 10, -1, -15, -5, 39, 19, -40, -1, 0, 39, -43, -7, -40, 15, -10, -4, -16, 5, -38, 56, 69, 44, -20, -33, 81, -19, -38, -6, 7, 7, -58, -32, 21, 49, -33, 48, -35, -1, 54, -10, -12, -15, -16, 16, -27, -7, -12, -13, -2, -4, -26, -54, 17, 45, 7, 34, -6, 29, -7, -5, -12, 34, 41, 59, -22, 29, -5, 16, -19, 22, -42, 12, -18, 13, 58, -56, -3, 3, 36, 19, -63, -17, -37, -12, -29, 12, -27, -36, 16, -33, -12, -3, 26, -12, 44, 49, 36, 37, 40, 15, -28, 12, -25, -13, -32, -43, 47, 37, -51, 38, 42, 56, 3, -46, 8, -46, 12, 51, 18, 4, -40, 66, 63, 45, -53, -95, 57, 61, -26, -4, 27, 34, 12, 36, -15, 32, -38, 1, -8, -25, -22, 24, -15, 19, -6, -27, 41, 17, 21, 13, 14, -4, -17, 31, -16, -32, 24, -22, -3, 31, -19, -21, 41, 8, -39, -8, 14, 22, -26, -3, 14, 13, -23, 38, 62, -42, -47, -16, 4, 33, -5, -37, 16, -17, 26, 11, 8, 6, -27, -3, -17, 9, 8, 35, 19, -14, 21, 36, 11, 43, 17, -21, -14, 16, -10, 48, -36, -27, 30, 50, 2, -37, -40, 38, -20, -2, 29, -58, -30, -77, -88, 15, -53, -58, 34, 8, -2, 34, -28, 2, 60, -20, -31, -17, 32, -29, -1, 42, 27, -11, 33, -22, -31, 21, 7, -40, 15, -1, 15, -14, -15, -1, -10, 6, -7, 51, 5, 0, -18, 55, 1, -14, 23, -11, 11, 37, -21, -64, -20, 12, 11, 43, 9, 41, 14, 26, 15, -47, -34, 0, 9, -7, -52, 8, -16, -28, 4, 32, 15, -13, -39, -29, -40, 21, 5, 34, -1, 28, -13, -13, 0, -15, -8, -16, -28, -12, -49, 12, -42, -61, -42, 11, -39, 1, 37, 0, 4, 4, -13, -45, -43, 6, 30, 62, 4, 7, 55, -6, -16, 27, -11, -14, -19, -16, -46, -8, -4, -19, -4, -15, 16, -35, -6, 27, 0, -18, 2, 28, 17, 38, -1, -1, 8, 14, 45, -13, -24, -2, 34, 40, 43, -36, -8, 53, 2, 21, 6, -51, -42, 29, -43, -2, -30, 12, 4, -20, 32, -50, -11, 34, 26, -29, 14, -47, -10, 11, -29, 25, 30, -34, -32, 19, 42, 1, -10, 7, 38, 29, 17, -11, -12, 20, -4, 48, 41, -41, -29, -6, -30, 24, -2, -11, 5, 10, 5, 7, -10, -5, 4, -27, -65, 36, 0, -33, -39, -12, -1, 17, 16, -40, -30, 2, -8, 25, 37, -9, 19, -23, 34, 12, -50, 7, 20, -6, -11, -7, 2, -3, -1, -9, -17, -40, 0, 1, -31, -43, -6, -27, 24, -29, 14, -13, -12, -1, 50, -24, 48, 29, 10, 2, 11, 14, -4, -13, 9, 10, 31, 11, -27, -5, 47, -17, 30, 25, 42, 26, 25, -4, -20, 15, 17, 1, 9, 54, 39, 46, -7, 1, 13, 14, 17, 55, 48, 56, 39, 35, 33, 39, 47, 46, -2, -3, 49, 4, -42, -14, -17, -5, 41, -25, 60, -6, -4, 59, 37, 23, 22, 27, 57, 22, 63, 16, 50, 28, 15, 40, 3, 5, 6, -39, 0, 9, 12, 5, -12, 0, 11, 20, -5, 21, 10, -1, -19, 11, 13, 28, -17, 33, -29, -9, -26, -15, 15, -10, 32, -38, 6, -10, -31, 14, 3, 36, -8, -4, -23, 15, -26, -29, 21, -16, 12, 0, -5, 32, 21, 53, -38, 4, 9, -20, 3, 0, 0, -6, 0, -3, 0, 0, -4, 0, 4, 4, 0, -4, 2, 0, 5, 0, -2, -3, 0, 0, 0, 0, 3, -1, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 4, -3, -2, 0, 5, 0, -2, 0, 2, 3, 0, 1, -1, -1, 0, 3, -1, 4, 0, -2, 0, -2, 0, 0, -3, 0, 0, -5, 0, 0, -2, 0, -2, -1, -1, 0, 0, 0, 0, 0, 2, 1, 0, 0, 3, 3, 0, 0, 0, -3, -3, 0, 0, -1, 0, 0, 0, -2, 0, 2, -5, -3, 1, 0, -1, 1, 4, -4, 0, 0, -3, 0, 0, 2, 0, -2, -1, 0, 0, 0, -1, 3, 0, 0, 0, 0, -1, 0, 0, 0, -1, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 1, -1, -2, 3, 0, -3, -5, 0, 0, 0, -1, 2, 0, 5, 2, 0, 0, 0, -4, 0, 0, 0, 0, 3, 0, 0, -3, -2, 0, -6, 0, 0, 0, 0, -5, -4, 0, 0, 0, 0, 1, 2, -2, 0, 2, -4, 0, -3, 4, -2, 0, -1, 0, 0, 0, 4, -6, 0, 0, 0, 0, -5, 19, 14, 8, 25, -1, 2, -33, -16, 10, 11, 2, 41, 1, 35, 25, -8, 31, 7, -28, 36, 34, 34, 2, -16, -30, 18, -34, -15, -31, -2, 4, -39, -38, -6, 36, 31, 6, -16, -57, -21, -8, -12, -5, -9, 3, 15, 16, -6, -48, -10, 23, -3, -20, -39, -46, 29, 22, 10, 6, 7, 41, 33, -14, 8, 25, -31, 2, -35, 1, -13, 5, -10, -24, -29, -19, 8, 32, -9, 10, 19, -49, -47, 16, 6, -8, -8, 8, 14, -34, 10, 12, 6, 52, 45, -10, -25, 11, 22, -24, -40, -38, -18, -10, -22, 1, 20, 25, -1, 19, 14, -26, -55, 46, -16, 28, -18, -6, 50, 36, -52, -55, 15, 49, 4, -56, 9, 49, 15, 12, 18, 7, -5, 6, -17, 18, -59, -51, -3, 26, 22, 16, -40, 12, 28, 25, 12, 24, 3, 14, 16, -4, -29, 32, 25, -47, -18, -9, 23, -3, -5, -33, 43, 13, 31, 1, -4, 24, -11, 28, 31, 14, -13, -20, 5, 25, 19, 34, -4, -8, 26, -47, 4, -16, 44, 30, 16, -34, 2, 28, 24, 48, 1, -13, 34, -11, -16, -10, 37, 28, -31, 31, 32, 2, 8, 3, 15, 40, 24, -27, -5, 27, 27, 10, 24, 41, -28, 23, 17, 28, 9, 2, 28, 18, 19, 8, -35, -38, -27, 20, 99, 14, -20, -8, 26, 60, -15, -40, 37, 2, -3, -13, -4, 8, -3, 3, 25, 36, -18, 13, -62, 19, 7, -13, -8, 25, -6, -21, -13, 18, 0, -24, -4, -13, 8, 44, 0, 7, 28, 43, 24, 22, 4, 17, -9, -2, 2, -1, 4, 2, -11, 21, 5, 17, 31, 40, -7, -22, -9, 28, -14, 24, -25, 13, -18, 52, -5, -1, 7, 7, -22, 18, 17, 48, -1, 37, 32, 15, 3, 49, 2, 48, 5, -52, -49, -43, -25, -70, 4, 5, 3, -21, -19, 34, -16, -46, 77, 75, 35, -14, -69, 60, 0, 59, 26, -24, 20, 19, -2, -22, 33, -40, 1, -19, 21, 56, -5, -15, -32, 10, 9, 5, -17, -34, 22, -5, -24, 30, 33, 3, 34, -21, 40, -30, -22, 4, 15, 63, -21, 24, 71, 4, -8, -10, -11, -69, -19, -3, -17, -27, -1, -23, 40, 28, 49, -22, 24, -19, -9, 43, 13, -22, -12, -55, -32, -7, 17, -12, 32, 17, -21, -7, -1, -27, 27, 9, -26, 28, -25, 38, 15, -23, -12, -31, -28, 22, 47, -1, -22, 31, -9, 23, 44, -35, -26, 19, -9, -19, -2, 45, 13, 29, -18, -23, 22, 64, 3, 4, -18, -10, -14, 21, -3, -10, -49, -53, -48, 25, -16, -1, -13, 10, -4, -22, -9, -38, -27, 2, -1, 7, -50, 34, 3, 7, 31, -12, -4, 48, -4, 32, 21, 25, 33, 15, -26, 14, -5, -27, 13, -31, 38, 29, 11, 30, 22, -11, -21, -33, -18, 7, 6, -24, -30, 2, 23, -29, 8, 19, 26, -1, -10, 26, 1, 22, 1, -30, 13, -2, 37, 4, -11, -15, -42, -13, -9, -3, -37, -9, -3, -3, -4, -66, -22, 35, -15, 50, 23, 37, 9, 17, -13, 26, 44, 26, 33, -29, 3, -10, 41, 5, -12, -20, -31, -13, -29, 19, 25, -23, 6, 59, 61, -11, -25, -25, -7, 15, 14, -11, 32, -21, -9, -22, -9, -6, -33, 30, 18, -17, -1, -3, -6, 26, 26, -1, 9, 26, 16, 36, -5, 11, -28, 2, -17, 34, 49, 7, 10, 24, -46, -36, 40, -23, 15, 9, -42, -21, -19, 41, 19, 8, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -21, -8, 29, 16, -50, 54, -19, -23, -29, -35, 25, 11, -33, -30, 8, -39, 21, 36, 25, -23, -2, -4, 43, 23, -28, -20, 12, -30, 17, -2, 30, -51, -19, 18, -22, 21, -1, 44, -28, 21, 2, 33, 44, -12, 20, -19, 15, 28, 22, -28, 33, 4, -16, -12, -22, 52, -5, -4, 35, 4, 4, 12, 24, 4, 11, -8, 30, 68, -51, 20, 13, 43, 3, -34, -18, 10, 23, 35, -2, 28, 60, -9, -15, -21, -7, -21, -53, -2, -18, -2, -20, -42, -7, 7, 25, -28, 35, 49, 3, 6, -35, -21, -36, -16, -28, 25, 27, -11, -15, -7, -54, -29, 19, 19, 13, -71, -10, 1, 26, 44, -50, -93, 40, 19, 23, 45, -3, -16, 52, 22, -22, 21, -23, 26, 12, 34, 16, -51, -55, 20, -40, -26, -66, 13, -16, -13, 24, -20, -2, 42, 20, 30, -8, 6, -6, 27, -12, -8, -29, 4, 15, -26, 2, -6, -3, 1, 9, 4, 22, 24, -13, -9, -10, 13, -24, -21, 45, 0, 50, -11, 56, 13, 17, 21, -10, -8, -11, 38, 3, -4, 24, -14, 41, -22, 8, -42, -10, 32, -42, -21, -4, -44, 8, -6, 31, -9, -4, 44, 21, 42, 20, 33, -4, 22, -5, 44, 13, 42, 41, -54, 29, 10, 7, 13, -2, 33, -48, 60, 40, 8, -9, -7, 39, -36, -20, 47, 31, 23, 62, 107, -18, 35, 32, -11, -27, 23, -20, 47, -5, -8, 34, 0, -26, -16, 46, -19, -6, 18, -16, 57, 7, -15, 27, -17, -39, 12, 12, 37, -28, -13, -34, 20, 61, 1, -96, -17, -28, 16, -46, 13, 29, -53, 39, -27, -7, -1, -39, 20, 4, -5, -6, -17, 27, 16, -61, 13, -10, 11, -10, -29, 18, -43, -60, 4, -45, 12, -16, -19, 26, 28, -2, 18, -79, 19, -19, 34, -7, 41, -9, -33, 10, -5, -16, -14, -26, -29, -64, -125, -67, 3, -21, -43, -38, -18, 30, -14, -46, -28, 49, -5, 59, -11, -62, -29, -36, 10, -6, 10, 25, -23, 7, -14, 18, 5, -1, 1, -44, 32, 41, 10, 31, -18, 18, 18, -48, 19, 19, 26, -27, -25, 29, 2, 44, -32, -53, -7, -39, -32, -44, -12, 26, -33, 8, 6, -7, -33, 3, 47, -30, 5, -1, -15, 46, -38, -62, -4, 40, 2, 13, 4, -2, 8, 29, 6, -29, 26, 43, -14, -25, 20, 29, -5, -48, 13, -8, -23, -10, 24, 28, 1, 31, -11, 36, 1, 39, 13, 41, -17, 11, 8, 16, 12, -13, 23, -17, 6, 12, -30, 27, 26, -9, -23, -20, -12, 4, -3, 12, -31, -44, 6, 8, 47, 9, -2, 33, 39, 39, -31, 12, -23, 26, -6, -28, -22, -38, -1, -7, -24, -4, 34, 38, 28, 0, 20, -39, -9, 50, -8, -14, -5, -14, 47, -10, -15, -24, 12, 38, -21, -31, 61, 30, -37, -20, -6, -26, -1, -8, 2, -35, 59, -14, 21, 19, -19, -42, -34, 21, 9, -2, 34, -34, -14, 47, -8, -2, -28, -2, 16, -18, -18, 15, -21, 49, 10, -21, -10, 4, 21, 20, 52, -30, -42, 10, -5, 28, -34, 5, -8, -13, -27, -26, 28, -19, -17, 41, -8, 49, 33, -2, 4, 16, 11, 19, 17, -22, -10, 46, 0, -6, 16, 4, 3, 7, -25, 9, -25, 26, -12, 3, 20, 7, -15, 47, 5, 11, -16, 28, 30, -21, -29, -3, -12, -35, -42, 9, 11, 28, -3, -35, 20, 27, 0, 19, -17, 8, -33, 8, 7, 19, -25, -5, -26, -24, 31, -22, 33, 28, 40, -6, -24, -2, -7, 24, 21, 17, -9, -9, -20, 10, -33, -24, -16, 11, 44, -18, 50, 47, 43, -20, -96, -11, -13, 8, 3, -32, 40, 45, -15, 14, 25, -18, -38, 37, -15, -14, 2, -7, 1, 42, 11, 27, 2, 7, 24, 34, 36, 63, -17, -32, 36, 14, -19, -43, 37, -10, -20, -38, 24, 5, 22, -15, 11, 49, 19, -4, 0, -11, -24, 18, 15, -22, 36, 12, -15, 6, 6, 33, -26, -13, -7, -1, 17, 19, -23, 7, -19, 30, 44, 15, -14, -24, -31, -23, 20, -14, -40, -48, 15, 37, 0, -15, 48, 58, 41, 3, 20, 38, -9, 18, -26, 6, 8, -51, 37, 36, -37, -5, -21, 15, 44, -53, -53, 6, 13, 66, 23, 13, 26, 1, 30, 59, 5, 45, -11, 9, -8, -3, -6, -30, -23, 2, 30, 7, 7, 37, -4, -6, 29, 39, -3, -11, -10, -6, 20, 6, 0, 22, 1, 37, -10, -6, -9, 12, 26, -6, 40, 11, 27, -36, -6, 52, 48, -18, -12, -40, 1, 33, -27, 37, 18, -20, 40, -21, -11, -27, -44, 4, 35, -15, 16, 11, 7, 25, 48, 27, 38, 40, -19, 31, 31, 14, -4, -27, 24, 12, -8, -23, -15, 37, -22, -12, 19, 1, -30, -20, -36, 9, -9, -57, -8, 9, -8, -17, 13, 35, -11, 52, -19, -5, 5, -30, 0, 25, 47, -15, 9, 22, 40, -16, -34, 18, -19, -25, -28, -7, 8, -34, 20, 23, 45, 25, 24, 39, 61, 40, 0, -44, -47, 46, 25, -32, 1, 9, 42, 11, -7, -16, 36, 40, -28, -19, -25, 42, 51, -17, -10, -4, -10, 20, 30, 20, -13, -14, 1, -4, -42, 3, 9, -24, -26, -6, 37, 47, 55, 19, -29, 4, -10, -35, 22, 8, -21, 8, 4, -20, -29, 71, 22, -37, -15, 15, 20, -40, -31, -20, -30, -11, 46, -26, -45, 24, 51, 40, 12, 26, -11, -5, -24, 59, 44, 6, 3, 50, 28, -49, 14, 21, 11, 5, -66, -30, -15, 13, 29, 7, 23, -27, -25, -18, -14, 9, 16, -12, 59, 36, 12, -29, -15, 28, -42, -32, -36, -5, -18, 17, -17, -31, 13, 14, 15, -1, -39, 7, -5, 39, 29, 33, -1, 57, 26, 1, 39, 14, 34, -28, 4, -19, 25, -12, 6, 14, -23, -32, -14, -9, 21, -18, 27, 10, 23, 29, 30, 29, 6, -19, 12, -6, -7, 2, 52, -27, 29, 32, 27, 14, 12, 23, -23, -2, -15, -39, -36, 16, -2, -24, -39, -1, -8, 3, 21, -13, 0, 22, 11, 9, -56, -1, 25, -54, -122, -10, 24, -13, -22, 11, 4, -3, 24, 11, 14, 26, 28, -1, -49, -8, 37, -1, -5, 43, -12, -52, 20, -22, 34, -56, 44, -9, 31, -6, 5, -29, -34, 13, 8, 15, -25, -12, -33, 30, -12, 14, -25, -30, 6, 21, -27, -3, 29, 10, -40, 26, 6, -6, -8, 21, 19, 45, 19, -10, 7, 27, 7, -49, 33, 57, 17, -17, 37, 28, -8, -28, 45, 23, -13, -26, -15, -1, 0, 17, -21, 25, 21, 18, 47, 2, -2, 41, 17, 5, -26, -22, 2, -30, 2, -7, -20, 26, -3, 0, -6, -19, -39, -16, -26, -4, -41, -9, -23, 18, -27, 19, 21, 10, -19, 40, 25, -1, -49, -28, 20, -10, -30, 16, -20, -11, 7, 34, -27, -36, 35, 0, -6, 10, -42, 24, -12, 4, -4, 26, 57, -1, -19,
    12, 37, 16, 34, -2, 26, -1, -9, 10, 19, -30, -22, 13, 44, -10, 5, 24, 8, 52, -7, -14, -44, 20, 16, 27, -36, -18, 26, 19, 3, -3, -33, -25, 7, 19, -12, 21, 66, -14, -9, -23, 14, 97, 9, -3, -23, -31, 66, 36, 2, -19, -28, 57, 22, -5, -14, 8, 29, 14, 34, -8, 26, 37, 12, -13, 5, -23, 2, 17, 32, -26, -18, 49, 38, 9, -23, 40, 25, -10, 26, 32, -18, 28, 21, 36, 14, 43, -1, -14, 10, -17, 9, 8, 24, -41, -43, -43, 39, 21, 12, -42, -27, 21, 39, -10, 11, 0, 31, 19, -27, 16, -5, -18, 26, 7, -7, -7, 9, 18, -12, -51, -18, -15, -45, 30, -20, -21, -8, 15, 22, 10, -14, -12, -26, 20, -2, 51, -7, -3, -1, -46, 1, 1, -58, -35, -34, -40, 10, 16, 10, -14, -20, 13, 20, 5, 11, 35, 21, 16, 7, -9, -6, 33, -7, 23, 0, -35, 38, 22, -9, 9, -7, 17, -8, 9, -31, 23, 16, 32, -33, 16, 7, -18, -18, 5, -28, -19, -23, 8, -22, -36, -32, 69, 8, -5, 11, -41, 37, 27, 2, -13, 19, 37, 25, 1, 13, -28, -2, -33, -19, 24, -11, 0, -11, 1, -24, -27, 28, -30, -4, 31, -5, 34, 47, -4, -7, 8, 27, 45, 13, -2, 29, -24, 2, -66, -18, -31, -46, -12, 23, 43, 29, 55, -35, -22, 46, 14, 8, -28, -14, -36, 16, -20, 16, 24, -2, 14, 17, 16, -8, -8, 8, -24, 18, -5, 4, 6, -69, 32, 5, -40, 3, -26, 30, -4, -19, 41, -45, 29, 19, -23, 8, 1, -20, -50, -39, 46, 17, -10, 19, 62, 64, 44, -43, -26, 8, -24, 22, -23, -13, -13, 17, -29, 12, 52, -32, -20, 10, -14, 2, 54, 32, 43, 29, -8, 3, 30, -1, 38, 22, 13, -20, -44, -32, -23, -23, 3, 33, 7, 43, 55, 9, -21, -27, -34, 28, 42, -34, -25, 11, 56, 38, 24, -1, 14, 21, 35, 1, -39, 28, -32, -34, -30, 2, 12, 9, -9, 40, -14, 27, 35, 26, 17, 37, -15, -33, 31, 14, 8, 22, 23, -20, -25, 37, -19, -42, -30, 34, -21, -13, -20, 2, 10, 33, -17, 11, -5, -16, -1, -35, 48, -2, 53, -37, -22, -5, -25, 50, -25, 17, -18, 1, -15, 7, 5, 18, 10, -11, 15, -7, -1, -15, -19, -16, 25, 37, -32, 16, 28, 39, -29, -26, -10, 35, -26, 44, -17, 6, 18, -20, -16, 31, -33, -5, 52, 15, 16, -36, 1, 8, 32, -16, -26, 30, 23, -11, 9, 44, 10, 26, 14, 10, 33, -19, 5, 22, 19, 39, 6, 50, 19, 50, 46, 52, 11, -13, 42, 2, 30, 1, -6, -13, -31, 19, 21, -11, 23, -9, -13, 6, 2, -32, 31, 19, -25, -22, -1, 44, 27, 28, -15, 3, 30, -11, -7, -25, 24, -15, 28, -17, -1, 30, -10, 35, 42, -2, 9, 0, -17, -35, -43, 21, -39, -41, -55, -51, -17, 8, -59, -12, 40, 37, -15, -64, -42, 33, 19, 10, -21, 5, 23, 8, 3, -19, -36, -38, 37, 27, -20, -46, -34, -12, 25, -26, -36, 3, 4, 22, -15, -28, 38, 20, 12, 8, 22, 34, 15, 4, -15, 34, 38, 46, 38, 25, 1, -30, -17, -36, -10, -10, -51, 19, -38, -11, -43, 39, 31, 24, -20, 33, -32, -15, 20, -18, -22, 42, 44, 9, 9, 21, 28, 7, -35, -14, 19, -12, 24, -33, 37, 55, 5, 5, 10, 5, 24, 43, 19, 39
  
  };

reg  signed [8:0] fc2_weights_re [0:639] = {

31, -63, 18, 28, -40, 19, -68, -88, -19, -31, 0, -62, 0, -28, -83, 52, 22, 14, 77, -86, 30, -37, -83, 70, -15, 72, 47, 62, -1, 47, -40, 28, -5, 79, -42, 26, -30, 81, -25, -74, -14, -59, -33, -19, 43, 16, 31, 3, -31, -64, 7, 56, 43, 80, 0, 27, -43, 27, -81, -10, 26, 42, 74, 54, 106, 74, -20, 8, -33, -31, 2, 59, -63, 74, 128, -28, 0, -33, -73, 8, 6, 7, -11, 4, 57, -39, 71, -23, 54, 74, 10, 52, -26, 23, 39, -5, 35, 4, -40, -4, 84, 44, 47, 102, 77, 31, 5, -93, 5, 1, -42, 57, 66, -93, 0, -85, -47, 0, 0, 35, 42, 12, 30, -89, -56, -13, -51, -6, 10, 69, 18, -61, -23, -120, -23, -47, 0, 60, 61, 25, 0, 23, -17, -77, -54, 84, 12, -75, -47, 82, 35, -62, 20, 42, -74, 17, 25, 83, 91, -65, -99, 74, 28, 98, 33, -35, 46, -47, 60, 53, 71, 80, -28, -54, -67, -12, 45, 5, 0, 36, 12, 93, 0, 4, -105, 36, -38, -83, -18, -48, 70, -15, -115, -89, -67, 46, -87, 4, 33, -23, -60, 45, -72, -17, 0, 30, -74, 80, 23, -12, 36, 41, 63, 73, 43, 23, -69, -5, -73, 59, 56, -65, -25, 57, -46, -30, 36, 15, 48, -53, 26, 50, 14, -17, 97, 68, 72, 65, -52, 41, -33, 68, -1, 63, -5, -4, 0, -79, -80, -88, -79, 28, 31, -29, -9, -86, -123, -47, 31, -97, 19, 47, -106, -112, 15, 60, 97, -23, 0, 82, 55, 47, -12, 4, -42, 50, -22, 73, 47, 13, 10, -38, 60, -66, -12, -45, -2, -86, -36, 82, 62, -78, 3, -88, -31, 10, 31, 53, -106, -70, -113, -27, 5, 16, -120, 32, 3, -21, -24, -1, 0, -92, -48, 32, 8, 11, -51, 47, -78, 49, 46, -34, -38, 17, -50, 44, -5, 70, -43, 79, 66, -42, 0, -27, 53, -3, 40, -20, 28, -17, 33, -54, -100, 57, -37, -126, -105, 88, 54, -22, -67, -67, -74, -52, -31, -85, 16, 72, -109, 75, -71, 16, -9, -35, 33, 74, 45, -72, -77, 73, 7, -58, -39, -43, 0, -57, 121, 70, 61, -37, 1, -137, 29, 1, 17, 47, 4, 19, -95, 57, 18, -29, 53, -18, -71, 72, 0, 72, 3, -9, -69, -68, 91, -43, 33, 26, -15, -50, 11, -48, -27, -67, -136, -1, -37, -75, -8, 22, -85, 35, 38, 44, -122, -20, 5, 74, 1, 27, -29, -51, 8, -149, -35, 52, -2, 52, -49, 4, 0, 83, 13, 67, 34, -79, 5, 17, -36, 78, 36, 169, 50, -86, -9, 79, -92, 6, -107, -67, 74, 43, 0, -6, 61, -20, 2, -46, 2, 70, -78, -91, -30, -4, 61, -81, -14, -32, -48, 20, -19, 39, -80, -32, -38, 72, -64, -52, 44, -1, 21, 48, 99, -55, -126, 55, 48, 73, 51, 66, 5, -60, 94, -24, 0, 42, -78, -44, 16, 48, 2, 15, 21, -78, 25, -25, -30, -56, -25, -38, -7, -25, 0, -90, -170, -86, 0, 43, 24, -148, -107, -64, 37, 76, -64, 33, -17, -47, 4, -17, -49, -2, 86, -12, 25, -45, -4, 20, 93, -4, 32, 51, -98, -90, -56, -42, -26, 15, 8, -7, -36, 4, -47, 38, -2, 13, 17, -23, 0, 25, -43, -9, -13, -9, -61, 5, 32, 45, 5, -147, -14, 40, 75, -79, -23, -61, -1, 60, 9, -86, 0, 41, 0, 82, -83, 69, -86, -16, -18, -18, -82, 55, 66, 74, -90, 61, 38, -39, -124, -24, -5, -2, -62, 85, -66, -46, -58, 14, 6, -187, -116, 15, -82, 4, -18, 7, 64, 22, 0, 17, -71, -45, 0, -152, -4, -18, 49, 89, -61, 61, 19, 37
};
