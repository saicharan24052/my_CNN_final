`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/17/2025 11:46:03 AM
// Design Name: 
// Module Name: add_conv2_modules
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module adder_28(
input logic clk,rst,
input logic signed [30:0] a,b,c,d,
output logic signed [32:0] sum
);

assign sum = a+b+c+d;


endmodule

module add_conv2_modules( // add 4 modules image1+img2+img3+img4 = output1
    input logic clk,rst,
    input logic signed [30:0] conv2_pre_final0 [0:120],
    input logic signed [30:0] conv2_pre_final1 [0:120],
    input logic signed [30:0] conv2_pre_final2 [0:120],
    input logic signed [30:0] conv2_pre_final3 [0:120],
    output logic signed [32:0] conv2_final_image [0:120]
    );
    
    
adder_28 mod28_0(clk,rst,conv2_pre_final0[0],conv2_pre_final1[0],conv2_pre_final2[0],conv2_pre_final3[0],conv2_final_image[0]);
    adder_28 mod28_1(clk,rst,conv2_pre_final0[1],conv2_pre_final1[1],conv2_pre_final2[1],conv2_pre_final3[1],conv2_final_image[1]);      
    adder_28 mod28_2(clk,rst,conv2_pre_final0[2],conv2_pre_final1[2],conv2_pre_final2[2],conv2_pre_final3[2],conv2_final_image[2]);      
    adder_28 mod28_3(clk,rst,conv2_pre_final0[3],conv2_pre_final1[3],conv2_pre_final2[3],conv2_pre_final3[3],conv2_final_image[3]);      
    adder_28 mod28_4(clk,rst,conv2_pre_final0[4],conv2_pre_final1[4],conv2_pre_final2[4],conv2_pre_final3[4],conv2_final_image[4]);      
    adder_28 mod28_5(clk,rst,conv2_pre_final0[5],conv2_pre_final1[5],conv2_pre_final2[5],conv2_pre_final3[5],conv2_final_image[5]);      
    adder_28 mod28_6(clk,rst,conv2_pre_final0[6],conv2_pre_final1[6],conv2_pre_final2[6],conv2_pre_final3[6],conv2_final_image[6]);      
    adder_28 mod28_7(clk,rst,conv2_pre_final0[7],conv2_pre_final1[7],conv2_pre_final2[7],conv2_pre_final3[7],conv2_final_image[7]);      
    adder_28 mod28_8(clk,rst,conv2_pre_final0[8],conv2_pre_final1[8],conv2_pre_final2[8],conv2_pre_final3[8],conv2_final_image[8]);      
    adder_28 mod28_9(clk,rst,conv2_pre_final0[9],conv2_pre_final1[9],conv2_pre_final2[9],conv2_pre_final3[9],conv2_final_image[9]);      
    adder_28 mod28_10(clk,rst,conv2_pre_final0[10],conv2_pre_final1[10],conv2_pre_final2[10],conv2_pre_final3[10],conv2_final_image[10]);
    adder_28 mod28_11(clk,rst,conv2_pre_final0[11],conv2_pre_final1[11],conv2_pre_final2[11],conv2_pre_final3[11],conv2_final_image[11]);
    adder_28 mod28_12(clk,rst,conv2_pre_final0[12],conv2_pre_final1[12],conv2_pre_final2[12],conv2_pre_final3[12],conv2_final_image[12]);
    adder_28 mod28_13(clk,rst,conv2_pre_final0[13],conv2_pre_final1[13],conv2_pre_final2[13],conv2_pre_final3[13],conv2_final_image[13]);
    adder_28 mod28_14(clk,rst,conv2_pre_final0[14],conv2_pre_final1[14],conv2_pre_final2[14],conv2_pre_final3[14],conv2_final_image[14]);
    adder_28 mod28_15(clk,rst,conv2_pre_final0[15],conv2_pre_final1[15],conv2_pre_final2[15],conv2_pre_final3[15],conv2_final_image[15]);
    adder_28 mod28_16(clk,rst,conv2_pre_final0[16],conv2_pre_final1[16],conv2_pre_final2[16],conv2_pre_final3[16],conv2_final_image[16]);
    adder_28 mod28_17(clk,rst,conv2_pre_final0[17],conv2_pre_final1[17],conv2_pre_final2[17],conv2_pre_final3[17],conv2_final_image[17]);
    adder_28 mod28_18(clk,rst,conv2_pre_final0[18],conv2_pre_final1[18],conv2_pre_final2[18],conv2_pre_final3[18],conv2_final_image[18]);
    adder_28 mod28_19(clk,rst,conv2_pre_final0[19],conv2_pre_final1[19],conv2_pre_final2[19],conv2_pre_final3[19],conv2_final_image[19]);
    adder_28 mod28_20(clk,rst,conv2_pre_final0[20],conv2_pre_final1[20],conv2_pre_final2[20],conv2_pre_final3[20],conv2_final_image[20]);
    adder_28 mod28_21(clk,rst,conv2_pre_final0[21],conv2_pre_final1[21],conv2_pre_final2[21],conv2_pre_final3[21],conv2_final_image[21]);
    adder_28 mod28_22(clk,rst,conv2_pre_final0[22],conv2_pre_final1[22],conv2_pre_final2[22],conv2_pre_final3[22],conv2_final_image[22]);
    adder_28 mod28_23(clk,rst,conv2_pre_final0[23],conv2_pre_final1[23],conv2_pre_final2[23],conv2_pre_final3[23],conv2_final_image[23]);
    adder_28 mod28_24(clk,rst,conv2_pre_final0[24],conv2_pre_final1[24],conv2_pre_final2[24],conv2_pre_final3[24],conv2_final_image[24]);
    adder_28 mod28_25(clk,rst,conv2_pre_final0[25],conv2_pre_final1[25],conv2_pre_final2[25],conv2_pre_final3[25],conv2_final_image[25]);
    adder_28 mod28_26(clk,rst,conv2_pre_final0[26],conv2_pre_final1[26],conv2_pre_final2[26],conv2_pre_final3[26],conv2_final_image[26]);
    adder_28 mod28_27(clk,rst,conv2_pre_final0[27],conv2_pre_final1[27],conv2_pre_final2[27],conv2_pre_final3[27],conv2_final_image[27]);
    adder_28 mod28_28(clk,rst,conv2_pre_final0[28],conv2_pre_final1[28],conv2_pre_final2[28],conv2_pre_final3[28],conv2_final_image[28]);
    adder_28 mod28_29(clk,rst,conv2_pre_final0[29],conv2_pre_final1[29],conv2_pre_final2[29],conv2_pre_final3[29],conv2_final_image[29]);
    adder_28 mod28_30(clk,rst,conv2_pre_final0[30],conv2_pre_final1[30],conv2_pre_final2[30],conv2_pre_final3[30],conv2_final_image[30]);
    adder_28 mod28_31(clk,rst,conv2_pre_final0[31],conv2_pre_final1[31],conv2_pre_final2[31],conv2_pre_final3[31],conv2_final_image[31]);
    adder_28 mod28_32(clk,rst,conv2_pre_final0[32],conv2_pre_final1[32],conv2_pre_final2[32],conv2_pre_final3[32],conv2_final_image[32]);
    adder_28 mod28_33(clk,rst,conv2_pre_final0[33],conv2_pre_final1[33],conv2_pre_final2[33],conv2_pre_final3[33],conv2_final_image[33]);
    adder_28 mod28_34(clk,rst,conv2_pre_final0[34],conv2_pre_final1[34],conv2_pre_final2[34],conv2_pre_final3[34],conv2_final_image[34]);
    adder_28 mod28_35(clk,rst,conv2_pre_final0[35],conv2_pre_final1[35],conv2_pre_final2[35],conv2_pre_final3[35],conv2_final_image[35]);
    adder_28 mod28_36(clk,rst,conv2_pre_final0[36],conv2_pre_final1[36],conv2_pre_final2[36],conv2_pre_final3[36],conv2_final_image[36]);
    adder_28 mod28_37(clk,rst,conv2_pre_final0[37],conv2_pre_final1[37],conv2_pre_final2[37],conv2_pre_final3[37],conv2_final_image[37]);
    adder_28 mod28_38(clk,rst,conv2_pre_final0[38],conv2_pre_final1[38],conv2_pre_final2[38],conv2_pre_final3[38],conv2_final_image[38]);
    adder_28 mod28_39(clk,rst,conv2_pre_final0[39],conv2_pre_final1[39],conv2_pre_final2[39],conv2_pre_final3[39],conv2_final_image[39]);
    adder_28 mod28_40(clk,rst,conv2_pre_final0[40],conv2_pre_final1[40],conv2_pre_final2[40],conv2_pre_final3[40],conv2_final_image[40]);
    adder_28 mod28_41(clk,rst,conv2_pre_final0[41],conv2_pre_final1[41],conv2_pre_final2[41],conv2_pre_final3[41],conv2_final_image[41]);
    adder_28 mod28_42(clk,rst,conv2_pre_final0[42],conv2_pre_final1[42],conv2_pre_final2[42],conv2_pre_final3[42],conv2_final_image[42]);
    adder_28 mod28_43(clk,rst,conv2_pre_final0[43],conv2_pre_final1[43],conv2_pre_final2[43],conv2_pre_final3[43],conv2_final_image[43]);
    adder_28 mod28_44(clk,rst,conv2_pre_final0[44],conv2_pre_final1[44],conv2_pre_final2[44],conv2_pre_final3[44],conv2_final_image[44]);
    adder_28 mod28_45(clk,rst,conv2_pre_final0[45],conv2_pre_final1[45],conv2_pre_final2[45],conv2_pre_final3[45],conv2_final_image[45]);
    adder_28 mod28_46(clk,rst,conv2_pre_final0[46],conv2_pre_final1[46],conv2_pre_final2[46],conv2_pre_final3[46],conv2_final_image[46]);
    adder_28 mod28_47(clk,rst,conv2_pre_final0[47],conv2_pre_final1[47],conv2_pre_final2[47],conv2_pre_final3[47],conv2_final_image[47]);
    adder_28 mod28_48(clk,rst,conv2_pre_final0[48],conv2_pre_final1[48],conv2_pre_final2[48],conv2_pre_final3[48],conv2_final_image[48]);
    adder_28 mod28_49(clk,rst,conv2_pre_final0[49],conv2_pre_final1[49],conv2_pre_final2[49],conv2_pre_final3[49],conv2_final_image[49]);
    adder_28 mod28_50(clk,rst,conv2_pre_final0[50],conv2_pre_final1[50],conv2_pre_final2[50],conv2_pre_final3[50],conv2_final_image[50]);
    adder_28 mod28_51(clk,rst,conv2_pre_final0[51],conv2_pre_final1[51],conv2_pre_final2[51],conv2_pre_final3[51],conv2_final_image[51]);
    adder_28 mod28_52(clk,rst,conv2_pre_final0[52],conv2_pre_final1[52],conv2_pre_final2[52],conv2_pre_final3[52],conv2_final_image[52]);
    adder_28 mod28_53(clk,rst,conv2_pre_final0[53],conv2_pre_final1[53],conv2_pre_final2[53],conv2_pre_final3[53],conv2_final_image[53]);
    adder_28 mod28_54(clk,rst,conv2_pre_final0[54],conv2_pre_final1[54],conv2_pre_final2[54],conv2_pre_final3[54],conv2_final_image[54]);
    adder_28 mod28_55(clk,rst,conv2_pre_final0[55],conv2_pre_final1[55],conv2_pre_final2[55],conv2_pre_final3[55],conv2_final_image[55]);
    adder_28 mod28_56(clk,rst,conv2_pre_final0[56],conv2_pre_final1[56],conv2_pre_final2[56],conv2_pre_final3[56],conv2_final_image[56]);
    adder_28 mod28_57(clk,rst,conv2_pre_final0[57],conv2_pre_final1[57],conv2_pre_final2[57],conv2_pre_final3[57],conv2_final_image[57]);
    adder_28 mod28_58(clk,rst,conv2_pre_final0[58],conv2_pre_final1[58],conv2_pre_final2[58],conv2_pre_final3[58],conv2_final_image[58]);
    adder_28 mod28_59(clk,rst,conv2_pre_final0[59],conv2_pre_final1[59],conv2_pre_final2[59],conv2_pre_final3[59],conv2_final_image[59]);
    adder_28 mod28_60(clk,rst,conv2_pre_final0[60],conv2_pre_final1[60],conv2_pre_final2[60],conv2_pre_final3[60],conv2_final_image[60]);
    adder_28 mod28_61(clk,rst,conv2_pre_final0[61],conv2_pre_final1[61],conv2_pre_final2[61],conv2_pre_final3[61],conv2_final_image[61]);
    adder_28 mod28_62(clk,rst,conv2_pre_final0[62],conv2_pre_final1[62],conv2_pre_final2[62],conv2_pre_final3[62],conv2_final_image[62]);
    adder_28 mod28_63(clk,rst,conv2_pre_final0[63],conv2_pre_final1[63],conv2_pre_final2[63],conv2_pre_final3[63],conv2_final_image[63]);
    adder_28 mod28_64(clk,rst,conv2_pre_final0[64],conv2_pre_final1[64],conv2_pre_final2[64],conv2_pre_final3[64],conv2_final_image[64]);
    adder_28 mod28_65(clk,rst,conv2_pre_final0[65],conv2_pre_final1[65],conv2_pre_final2[65],conv2_pre_final3[65],conv2_final_image[65]);
    adder_28 mod28_66(clk,rst,conv2_pre_final0[66],conv2_pre_final1[66],conv2_pre_final2[66],conv2_pre_final3[66],conv2_final_image[66]);
    adder_28 mod28_67(clk,rst,conv2_pre_final0[67],conv2_pre_final1[67],conv2_pre_final2[67],conv2_pre_final3[67],conv2_final_image[67]);
    adder_28 mod28_68(clk,rst,conv2_pre_final0[68],conv2_pre_final1[68],conv2_pre_final2[68],conv2_pre_final3[68],conv2_final_image[68]);
    adder_28 mod28_69(clk,rst,conv2_pre_final0[69],conv2_pre_final1[69],conv2_pre_final2[69],conv2_pre_final3[69],conv2_final_image[69]);
    adder_28 mod28_70(clk,rst,conv2_pre_final0[70],conv2_pre_final1[70],conv2_pre_final2[70],conv2_pre_final3[70],conv2_final_image[70]);
    adder_28 mod28_71(clk,rst,conv2_pre_final0[71],conv2_pre_final1[71],conv2_pre_final2[71],conv2_pre_final3[71],conv2_final_image[71]);
    adder_28 mod28_72(clk,rst,conv2_pre_final0[72],conv2_pre_final1[72],conv2_pre_final2[72],conv2_pre_final3[72],conv2_final_image[72]);
    adder_28 mod28_73(clk,rst,conv2_pre_final0[73],conv2_pre_final1[73],conv2_pre_final2[73],conv2_pre_final3[73],conv2_final_image[73]);
    adder_28 mod28_74(clk,rst,conv2_pre_final0[74],conv2_pre_final1[74],conv2_pre_final2[74],conv2_pre_final3[74],conv2_final_image[74]);
    adder_28 mod28_75(clk,rst,conv2_pre_final0[75],conv2_pre_final1[75],conv2_pre_final2[75],conv2_pre_final3[75],conv2_final_image[75]);
    adder_28 mod28_76(clk,rst,conv2_pre_final0[76],conv2_pre_final1[76],conv2_pre_final2[76],conv2_pre_final3[76],conv2_final_image[76]);
    adder_28 mod28_77(clk,rst,conv2_pre_final0[77],conv2_pre_final1[77],conv2_pre_final2[77],conv2_pre_final3[77],conv2_final_image[77]);
    adder_28 mod28_78(clk,rst,conv2_pre_final0[78],conv2_pre_final1[78],conv2_pre_final2[78],conv2_pre_final3[78],conv2_final_image[78]);
    adder_28 mod28_79(clk,rst,conv2_pre_final0[79],conv2_pre_final1[79],conv2_pre_final2[79],conv2_pre_final3[79],conv2_final_image[79]);
    adder_28 mod28_80(clk,rst,conv2_pre_final0[80],conv2_pre_final1[80],conv2_pre_final2[80],conv2_pre_final3[80],conv2_final_image[80]);
    adder_28 mod28_81(clk,rst,conv2_pre_final0[81],conv2_pre_final1[81],conv2_pre_final2[81],conv2_pre_final3[81],conv2_final_image[81]);
    adder_28 mod28_82(clk,rst,conv2_pre_final0[82],conv2_pre_final1[82],conv2_pre_final2[82],conv2_pre_final3[82],conv2_final_image[82]);
    adder_28 mod28_83(clk,rst,conv2_pre_final0[83],conv2_pre_final1[83],conv2_pre_final2[83],conv2_pre_final3[83],conv2_final_image[83]);
    adder_28 mod28_84(clk,rst,conv2_pre_final0[84],conv2_pre_final1[84],conv2_pre_final2[84],conv2_pre_final3[84],conv2_final_image[84]);
    adder_28 mod28_85(clk,rst,conv2_pre_final0[85],conv2_pre_final1[85],conv2_pre_final2[85],conv2_pre_final3[85],conv2_final_image[85]);
    adder_28 mod28_86(clk,rst,conv2_pre_final0[86],conv2_pre_final1[86],conv2_pre_final2[86],conv2_pre_final3[86],conv2_final_image[86]);
    adder_28 mod28_87(clk,rst,conv2_pre_final0[87],conv2_pre_final1[87],conv2_pre_final2[87],conv2_pre_final3[87],conv2_final_image[87]);
    adder_28 mod28_88(clk,rst,conv2_pre_final0[88],conv2_pre_final1[88],conv2_pre_final2[88],conv2_pre_final3[88],conv2_final_image[88]);
    adder_28 mod28_89(clk,rst,conv2_pre_final0[89],conv2_pre_final1[89],conv2_pre_final2[89],conv2_pre_final3[89],conv2_final_image[89]);
    adder_28 mod28_90(clk,rst,conv2_pre_final0[90],conv2_pre_final1[90],conv2_pre_final2[90],conv2_pre_final3[90],conv2_final_image[90]);
    adder_28 mod28_91(clk,rst,conv2_pre_final0[91],conv2_pre_final1[91],conv2_pre_final2[91],conv2_pre_final3[91],conv2_final_image[91]);
    adder_28 mod28_92(clk,rst,conv2_pre_final0[92],conv2_pre_final1[92],conv2_pre_final2[92],conv2_pre_final3[92],conv2_final_image[92]);
    adder_28 mod28_93(clk,rst,conv2_pre_final0[93],conv2_pre_final1[93],conv2_pre_final2[93],conv2_pre_final3[93],conv2_final_image[93]);
    adder_28 mod28_94(clk,rst,conv2_pre_final0[94],conv2_pre_final1[94],conv2_pre_final2[94],conv2_pre_final3[94],conv2_final_image[94]);
    adder_28 mod28_95(clk,rst,conv2_pre_final0[95],conv2_pre_final1[95],conv2_pre_final2[95],conv2_pre_final3[95],conv2_final_image[95]);
    adder_28 mod28_96(clk,rst,conv2_pre_final0[96],conv2_pre_final1[96],conv2_pre_final2[96],conv2_pre_final3[96],conv2_final_image[96]);
    adder_28 mod28_97(clk,rst,conv2_pre_final0[97],conv2_pre_final1[97],conv2_pre_final2[97],conv2_pre_final3[97],conv2_final_image[97]);
    adder_28 mod28_98(clk,rst,conv2_pre_final0[98],conv2_pre_final1[98],conv2_pre_final2[98],conv2_pre_final3[98],conv2_final_image[98]);
    adder_28 mod28_99(clk,rst,conv2_pre_final0[99],conv2_pre_final1[99],conv2_pre_final2[99],conv2_pre_final3[99],conv2_final_image[99]);
    adder_28 mod28_100(clk,rst,conv2_pre_final0[100],conv2_pre_final1[100],conv2_pre_final2[100],conv2_pre_final3[100],conv2_final_image[100]);
    adder_28 mod28_101(clk,rst,conv2_pre_final0[101],conv2_pre_final1[101],conv2_pre_final2[101],conv2_pre_final3[101],conv2_final_image[101]);
    adder_28 mod28_102(clk,rst,conv2_pre_final0[102],conv2_pre_final1[102],conv2_pre_final2[102],conv2_pre_final3[102],conv2_final_image[102]);
    adder_28 mod28_103(clk,rst,conv2_pre_final0[103],conv2_pre_final1[103],conv2_pre_final2[103],conv2_pre_final3[103],conv2_final_image[103]);
    adder_28 mod28_104(clk,rst,conv2_pre_final0[104],conv2_pre_final1[104],conv2_pre_final2[104],conv2_pre_final3[104],conv2_final_image[104]);
    adder_28 mod28_105(clk,rst,conv2_pre_final0[105],conv2_pre_final1[105],conv2_pre_final2[105],conv2_pre_final3[105],conv2_final_image[105]);
    adder_28 mod28_106(clk,rst,conv2_pre_final0[106],conv2_pre_final1[106],conv2_pre_final2[106],conv2_pre_final3[106],conv2_final_image[106]);
    adder_28 mod28_107(clk,rst,conv2_pre_final0[107],conv2_pre_final1[107],conv2_pre_final2[107],conv2_pre_final3[107],conv2_final_image[107]);
    adder_28 mod28_108(clk,rst,conv2_pre_final0[108],conv2_pre_final1[108],conv2_pre_final2[108],conv2_pre_final3[108],conv2_final_image[108]);
    adder_28 mod28_109(clk,rst,conv2_pre_final0[109],conv2_pre_final1[109],conv2_pre_final2[109],conv2_pre_final3[109],conv2_final_image[109]);
    adder_28 mod28_110(clk,rst,conv2_pre_final0[110],conv2_pre_final1[110],conv2_pre_final2[110],conv2_pre_final3[110],conv2_final_image[110]);
    adder_28 mod28_111(clk,rst,conv2_pre_final0[111],conv2_pre_final1[111],conv2_pre_final2[111],conv2_pre_final3[111],conv2_final_image[111]);
    adder_28 mod28_112(clk,rst,conv2_pre_final0[112],conv2_pre_final1[112],conv2_pre_final2[112],conv2_pre_final3[112],conv2_final_image[112]);
    adder_28 mod28_113(clk,rst,conv2_pre_final0[113],conv2_pre_final1[113],conv2_pre_final2[113],conv2_pre_final3[113],conv2_final_image[113]);
    adder_28 mod28_114(clk,rst,conv2_pre_final0[114],conv2_pre_final1[114],conv2_pre_final2[114],conv2_pre_final3[114],conv2_final_image[114]);
    adder_28 mod28_115(clk,rst,conv2_pre_final0[115],conv2_pre_final1[115],conv2_pre_final2[115],conv2_pre_final3[115],conv2_final_image[115]);
    adder_28 mod28_116(clk,rst,conv2_pre_final0[116],conv2_pre_final1[116],conv2_pre_final2[116],conv2_pre_final3[116],conv2_final_image[116]);
    adder_28 mod28_117(clk,rst,conv2_pre_final0[117],conv2_pre_final1[117],conv2_pre_final2[117],conv2_pre_final3[117],conv2_final_image[117]);
    adder_28 mod28_118(clk,rst,conv2_pre_final0[118],conv2_pre_final1[118],conv2_pre_final2[118],conv2_pre_final3[118],conv2_final_image[118]);
    adder_28 mod28_119(clk,rst,conv2_pre_final0[119],conv2_pre_final1[119],conv2_pre_final2[119],conv2_pre_final3[119],conv2_final_image[119]);
    adder_28 mod28_120(clk,rst,conv2_pre_final0[120],conv2_pre_final1[120],conv2_pre_final2[120],conv2_pre_final3[120],conv2_final_image[120]);
    
    
    
    
    
    
    
    
    
    
    
endmodule
