`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/11/2025 03:13:16 PM
// Design Name: 
// Module Name: CNN_conv2_final_mod
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module adder_24bit ( // with sign
input logic signed [26:0]aa,bb,cc,dd,ee,ff,gg,hh,hhi,
output logic signed [30:0] sum2 //signed
);

assign sum2 = aa+bb+cc+dd+ee+ff+gg+hh+hhi; // add all without sign bit
endmodule


module mul_20x8bit(
input logic signed [19:0]aal, // 8bit a without signed and 8 bit 256
input logic signed [7:0]bbl, // max number after mul with 256 is 63(6bit)7 bit with sign
output logic signed [26:0] multi_out2
);

assign multi_out2 = aal*bbl; // multiply all without sign bit al[7:0]*bl[5:0]
endmodule


 module CNN_conv2_final_mod(
input logic clk,rst,
input logic signed [19:0] image2[0:168], // unsigned
input logic signed [7:0]filter_2[0:8], // signed(max:63) kernel_1_re[4]3][3]: kernel_1_re[0][x][y],kernel_1_re[1][x][y], . kernel_1_re[3][x][y], round off 3 decimal points
output logic signed [30:0] conv2_out [0:120] // signed
);
 logic signed [26:0] mul2_out [0:362][0:12]; // signed

mul_20x8bit m2_0 (image2[0],filter_2[0],mul2_out[0][0]);
mul_20x8bit m2_1 (image2[1],filter_2[1],mul2_out[0][1]);
mul_20x8bit m2_2 (image2[2],filter_2[2],mul2_out[0][2]);
mul_20x8bit m2_3 (image2[13],filter_2[3],mul2_out[1][0]);
mul_20x8bit m2_4 (image2[14],filter_2[4],mul2_out[1][1]);
mul_20x8bit m2_5 (image2[15],filter_2[5],mul2_out[1][2]);
mul_20x8bit m2_6 (image2[26],filter_2[6],mul2_out[2][0]);
mul_20x8bit m2_7 (image2[27],filter_2[7],mul2_out[2][1]);
mul_20x8bit m2_8 (image2[28],filter_2[8],mul2_out[2][2]);

adder_24bit ad2_0 (mul2_out[0][0],mul2_out[0][1],mul2_out[0][2],mul2_out[1][0],mul2_out[1][1],mul2_out[1][2],mul2_out[2][0],mul2_out[2][1],mul2_out[2][2],conv2_out[0]);



mul_20x8bit m2_9 (image2[1],filter_2[0],mul2_out[3][0]);
mul_20x8bit m2_10 (image2[2],filter_2[1],mul2_out[3][1]);
mul_20x8bit m2_11 (image2[3],filter_2[2],mul2_out[3][2]);
mul_20x8bit m2_12 (image2[14],filter_2[3],mul2_out[4][0]);
mul_20x8bit m2_13 (image2[15],filter_2[4],mul2_out[4][1]);
mul_20x8bit m2_14 (image2[16],filter_2[5],mul2_out[4][2]);
mul_20x8bit m2_15 (image2[27],filter_2[6],mul2_out[5][0]);
mul_20x8bit m2_16 (image2[28],filter_2[7],mul2_out[5][1]);
mul_20x8bit m2_17 (image2[29],filter_2[8],mul2_out[5][2]);

adder_24bit ad2_1 (mul2_out[3][0],mul2_out[3][1],mul2_out[3][2],mul2_out[4][0],mul2_out[4][1],mul2_out[4][2],mul2_out[5][0],mul2_out[5][1],mul2_out[5][2],conv2_out[1]);



mul_20x8bit m2_18 (image2[2],filter_2[0],mul2_out[6][0]);
mul_20x8bit m2_19 (image2[3],filter_2[1],mul2_out[6][1]);
mul_20x8bit m2_20 (image2[4],filter_2[2],mul2_out[6][2]);
mul_20x8bit m2_21 (image2[15],filter_2[3],mul2_out[7][0]);
mul_20x8bit m2_22 (image2[16],filter_2[4],mul2_out[7][1]);
mul_20x8bit m2_23 (image2[17],filter_2[5],mul2_out[7][2]);
mul_20x8bit m2_24 (image2[28],filter_2[6],mul2_out[8][0]);
mul_20x8bit m2_25 (image2[29],filter_2[7],mul2_out[8][1]);
mul_20x8bit m2_26 (image2[30],filter_2[8],mul2_out[8][2]);

adder_24bit ad2_2 (mul2_out[6][0],mul2_out[6][1],mul2_out[6][2],mul2_out[7][0],mul2_out[7][1],mul2_out[7][2],mul2_out[8][0],mul2_out[8][1],mul2_out[8][2],conv2_out[2]);



mul_20x8bit m2_27 (image2[3],filter_2[0],mul2_out[9][0]);
mul_20x8bit m2_28 (image2[4],filter_2[1],mul2_out[9][1]);
mul_20x8bit m2_29 (image2[5],filter_2[2],mul2_out[9][2]);
mul_20x8bit m2_30 (image2[16],filter_2[3],mul2_out[10][0]);
mul_20x8bit m2_31 (image2[17],filter_2[4],mul2_out[10][1]);
mul_20x8bit m2_32 (image2[18],filter_2[5],mul2_out[10][2]);
mul_20x8bit m2_33 (image2[29],filter_2[6],mul2_out[11][0]);
mul_20x8bit m2_34 (image2[30],filter_2[7],mul2_out[11][1]);
mul_20x8bit m2_35 (image2[31],filter_2[8],mul2_out[11][2]);

adder_24bit ad2_3 (mul2_out[9][0],mul2_out[9][1],mul2_out[9][2],mul2_out[10][0],mul2_out[10][1],mul2_out[10][2],mul2_out[11][0],mul2_out[11][1],mul2_out[11][2],conv2_out[3]);



mul_20x8bit m2_36 (image2[4],filter_2[0],mul2_out[12][0]);
mul_20x8bit m2_37 (image2[5],filter_2[1],mul2_out[12][1]);
mul_20x8bit m2_38 (image2[6],filter_2[2],mul2_out[12][2]);
mul_20x8bit m2_39 (image2[17],filter_2[3],mul2_out[13][0]);
mul_20x8bit m2_40 (image2[18],filter_2[4],mul2_out[13][1]);
mul_20x8bit m2_41 (image2[19],filter_2[5],mul2_out[13][2]);
mul_20x8bit m2_42 (image2[30],filter_2[6],mul2_out[14][0]);
mul_20x8bit m2_43 (image2[31],filter_2[7],mul2_out[14][1]);
mul_20x8bit m2_44 (image2[32],filter_2[8],mul2_out[14][2]);

adder_24bit ad2_4 (mul2_out[12][0],mul2_out[12][1],mul2_out[12][2],mul2_out[13][0],mul2_out[13][1],mul2_out[13][2],mul2_out[14][0],mul2_out[14][1],mul2_out[14][2],conv2_out[4]);



mul_20x8bit m2_45 (image2[5],filter_2[0],mul2_out[15][0]);
mul_20x8bit m2_46 (image2[6],filter_2[1],mul2_out[15][1]);
mul_20x8bit m2_47 (image2[7],filter_2[2],mul2_out[15][2]);
mul_20x8bit m2_48 (image2[18],filter_2[3],mul2_out[16][0]);
mul_20x8bit m2_49 (image2[19],filter_2[4],mul2_out[16][1]);
mul_20x8bit m2_50 (image2[20],filter_2[5],mul2_out[16][2]);
mul_20x8bit m2_51 (image2[31],filter_2[6],mul2_out[17][0]);
mul_20x8bit m2_52 (image2[32],filter_2[7],mul2_out[17][1]);
mul_20x8bit m2_53 (image2[33],filter_2[8],mul2_out[17][2]);

adder_24bit ad2_5 (mul2_out[15][0],mul2_out[15][1],mul2_out[15][2],mul2_out[16][0],mul2_out[16][1],mul2_out[16][2],mul2_out[17][0],mul2_out[17][1],mul2_out[17][2],conv2_out[5]);



mul_20x8bit m2_54 (image2[6],filter_2[0],mul2_out[18][0]);
mul_20x8bit m2_55 (image2[7],filter_2[1],mul2_out[18][1]);
mul_20x8bit m2_56 (image2[8],filter_2[2],mul2_out[18][2]);
mul_20x8bit m2_57 (image2[19],filter_2[3],mul2_out[19][0]);
mul_20x8bit m2_58 (image2[20],filter_2[4],mul2_out[19][1]);
mul_20x8bit m2_59 (image2[21],filter_2[5],mul2_out[19][2]);
mul_20x8bit m2_60 (image2[32],filter_2[6],mul2_out[20][0]);
mul_20x8bit m2_61 (image2[33],filter_2[7],mul2_out[20][1]);
mul_20x8bit m2_62 (image2[34],filter_2[8],mul2_out[20][2]);

adder_24bit ad2_6 (mul2_out[18][0],mul2_out[18][1],mul2_out[18][2],mul2_out[19][0],mul2_out[19][1],mul2_out[19][2],mul2_out[20][0],mul2_out[20][1],mul2_out[20][2],conv2_out[6]);



mul_20x8bit m2_63 (image2[7],filter_2[0],mul2_out[21][0]);
mul_20x8bit m2_64 (image2[8],filter_2[1],mul2_out[21][1]);
mul_20x8bit m2_65 (image2[9],filter_2[2],mul2_out[21][2]);
mul_20x8bit m2_66 (image2[20],filter_2[3],mul2_out[22][0]);
mul_20x8bit m2_67 (image2[21],filter_2[4],mul2_out[22][1]);
mul_20x8bit m2_68 (image2[22],filter_2[5],mul2_out[22][2]);
mul_20x8bit m2_69 (image2[33],filter_2[6],mul2_out[23][0]);
mul_20x8bit m2_70 (image2[34],filter_2[7],mul2_out[23][1]);
mul_20x8bit m2_71 (image2[35],filter_2[8],mul2_out[23][2]);

adder_24bit ad2_7 (mul2_out[21][0],mul2_out[21][1],mul2_out[21][2],mul2_out[22][0],mul2_out[22][1],mul2_out[22][2],mul2_out[23][0],mul2_out[23][1],mul2_out[23][2],conv2_out[7]);



mul_20x8bit m2_72 (image2[8],filter_2[0],mul2_out[24][0]);
mul_20x8bit m2_73 (image2[9],filter_2[1],mul2_out[24][1]);
mul_20x8bit m2_74 (image2[10],filter_2[2],mul2_out[24][2]);
mul_20x8bit m2_75 (image2[21],filter_2[3],mul2_out[25][0]);
mul_20x8bit m2_76 (image2[22],filter_2[4],mul2_out[25][1]);
mul_20x8bit m2_77 (image2[23],filter_2[5],mul2_out[25][2]);
mul_20x8bit m2_78 (image2[34],filter_2[6],mul2_out[26][0]);
mul_20x8bit m2_79 (image2[35],filter_2[7],mul2_out[26][1]);
mul_20x8bit m2_80 (image2[36],filter_2[8],mul2_out[26][2]);

adder_24bit ad2_8 (mul2_out[24][0],mul2_out[24][1],mul2_out[24][2],mul2_out[25][0],mul2_out[25][1],mul2_out[25][2],mul2_out[26][0],mul2_out[26][1],mul2_out[26][2],conv2_out[8]);



mul_20x8bit m2_81 (image2[9],filter_2[0],mul2_out[27][0]);
mul_20x8bit m2_82 (image2[10],filter_2[1],mul2_out[27][1]);
mul_20x8bit m2_83 (image2[11],filter_2[2],mul2_out[27][2]);
mul_20x8bit m2_84 (image2[22],filter_2[3],mul2_out[28][0]);
mul_20x8bit m2_85 (image2[23],filter_2[4],mul2_out[28][1]);
mul_20x8bit m2_86 (image2[24],filter_2[5],mul2_out[28][2]);
mul_20x8bit m2_87 (image2[35],filter_2[6],mul2_out[29][0]);
mul_20x8bit m2_88 (image2[36],filter_2[7],mul2_out[29][1]);
mul_20x8bit m2_89 (image2[37],filter_2[8],mul2_out[29][2]);

adder_24bit ad2_9 (mul2_out[27][0],mul2_out[27][1],mul2_out[27][2],mul2_out[28][0],mul2_out[28][1],mul2_out[28][2],mul2_out[29][0],mul2_out[29][1],mul2_out[29][2],conv2_out[9]);



mul_20x8bit m2_90 (image2[10],filter_2[0],mul2_out[30][0]);
mul_20x8bit m2_91 (image2[11],filter_2[1],mul2_out[30][1]);
mul_20x8bit m2_92 (image2[12],filter_2[2],mul2_out[30][2]);
mul_20x8bit m2_93 (image2[23],filter_2[3],mul2_out[31][0]);
mul_20x8bit m2_94 (image2[24],filter_2[4],mul2_out[31][1]);
mul_20x8bit m2_95 (image2[25],filter_2[5],mul2_out[31][2]);
mul_20x8bit m2_96 (image2[36],filter_2[6],mul2_out[32][0]);
mul_20x8bit m2_97 (image2[37],filter_2[7],mul2_out[32][1]);
mul_20x8bit m2_98 (image2[38],filter_2[8],mul2_out[32][2]);

adder_24bit ad2_10 (mul2_out[30][0],mul2_out[30][1],mul2_out[30][2],mul2_out[31][0],mul2_out[31][1],mul2_out[31][2],mul2_out[32][0],mul2_out[32][1],mul2_out[32][2],conv2_out[10]);



mul_20x8bit m2_99 (image2[13],filter_2[0],mul2_out[33][1]);
mul_20x8bit m2_100 (image2[14],filter_2[1],mul2_out[33][2]);
mul_20x8bit m2_101 (image2[15],filter_2[2],mul2_out[33][3]);
mul_20x8bit m2_102 (image2[26],filter_2[3],mul2_out[34][1]);
mul_20x8bit m2_103 (image2[27],filter_2[4],mul2_out[34][2]);
mul_20x8bit m2_104 (image2[28],filter_2[5],mul2_out[34][3]);
mul_20x8bit m2_105 (image2[39],filter_2[6],mul2_out[35][1]);
mul_20x8bit m2_106 (image2[40],filter_2[7],mul2_out[35][2]);
mul_20x8bit m2_107 (image2[41],filter_2[8],mul2_out[35][3]);

adder_24bit ad2_11 (mul2_out[33][1],mul2_out[33][2],mul2_out[33][3],mul2_out[34][1],mul2_out[34][2],mul2_out[34][3],mul2_out[35][1],mul2_out[35][2],mul2_out[35][3],conv2_out[11]);



mul_20x8bit m2_108 (image2[14],filter_2[0],mul2_out[36][1]);
mul_20x8bit m2_109 (image2[15],filter_2[1],mul2_out[36][2]);
mul_20x8bit m2_110 (image2[16],filter_2[2],mul2_out[36][3]);
mul_20x8bit m2_111 (image2[27],filter_2[3],mul2_out[37][1]);
mul_20x8bit m2_112 (image2[28],filter_2[4],mul2_out[37][2]);
mul_20x8bit m2_113 (image2[29],filter_2[5],mul2_out[37][3]);
mul_20x8bit m2_114 (image2[40],filter_2[6],mul2_out[38][1]);
mul_20x8bit m2_115 (image2[41],filter_2[7],mul2_out[38][2]);
mul_20x8bit m2_116 (image2[42],filter_2[8],mul2_out[38][3]);

adder_24bit ad2_12 (mul2_out[36][1],mul2_out[36][2],mul2_out[36][3],mul2_out[37][1],mul2_out[37][2],mul2_out[37][3],mul2_out[38][1],mul2_out[38][2],mul2_out[38][3],conv2_out[12]);



mul_20x8bit m2_117 (image2[15],filter_2[0],mul2_out[39][1]);
mul_20x8bit m2_118 (image2[16],filter_2[1],mul2_out[39][2]);
mul_20x8bit m2_119 (image2[17],filter_2[2],mul2_out[39][3]);
mul_20x8bit m2_120 (image2[28],filter_2[3],mul2_out[40][1]);
mul_20x8bit m2_121 (image2[29],filter_2[4],mul2_out[40][2]);
mul_20x8bit m2_122 (image2[30],filter_2[5],mul2_out[40][3]);
mul_20x8bit m2_123 (image2[41],filter_2[6],mul2_out[41][1]);
mul_20x8bit m2_124 (image2[42],filter_2[7],mul2_out[41][2]);
mul_20x8bit m2_125 (image2[43],filter_2[8],mul2_out[41][3]);

adder_24bit ad2_13 (mul2_out[39][1],mul2_out[39][2],mul2_out[39][3],mul2_out[40][1],mul2_out[40][2],mul2_out[40][3],mul2_out[41][1],mul2_out[41][2],mul2_out[41][3],conv2_out[13]);



mul_20x8bit m2_126 (image2[16],filter_2[0],mul2_out[42][1]);
mul_20x8bit m2_127 (image2[17],filter_2[1],mul2_out[42][2]);
mul_20x8bit m2_128 (image2[18],filter_2[2],mul2_out[42][3]);
mul_20x8bit m2_129 (image2[29],filter_2[3],mul2_out[43][1]);
mul_20x8bit m2_130 (image2[30],filter_2[4],mul2_out[43][2]);
mul_20x8bit m2_131 (image2[31],filter_2[5],mul2_out[43][3]);
mul_20x8bit m2_132 (image2[42],filter_2[6],mul2_out[44][1]);
mul_20x8bit m2_133 (image2[43],filter_2[7],mul2_out[44][2]);
mul_20x8bit m2_134 (image2[44],filter_2[8],mul2_out[44][3]);

adder_24bit ad2_14 (mul2_out[42][1],mul2_out[42][2],mul2_out[42][3],mul2_out[43][1],mul2_out[43][2],mul2_out[43][3],mul2_out[44][1],mul2_out[44][2],mul2_out[44][3],conv2_out[14]);



mul_20x8bit m2_135 (image2[17],filter_2[0],mul2_out[45][1]);
mul_20x8bit m2_136 (image2[18],filter_2[1],mul2_out[45][2]);
mul_20x8bit m2_137 (image2[19],filter_2[2],mul2_out[45][3]);
mul_20x8bit m2_138 (image2[30],filter_2[3],mul2_out[46][1]);
mul_20x8bit m2_139 (image2[31],filter_2[4],mul2_out[46][2]);
mul_20x8bit m2_140 (image2[32],filter_2[5],mul2_out[46][3]);
mul_20x8bit m2_141 (image2[43],filter_2[6],mul2_out[47][1]);
mul_20x8bit m2_142 (image2[44],filter_2[7],mul2_out[47][2]);
mul_20x8bit m2_143 (image2[45],filter_2[8],mul2_out[47][3]);

adder_24bit ad2_15 (mul2_out[45][1],mul2_out[45][2],mul2_out[45][3],mul2_out[46][1],mul2_out[46][2],mul2_out[46][3],mul2_out[47][1],mul2_out[47][2],mul2_out[47][3],conv2_out[15]);



mul_20x8bit m2_144 (image2[18],filter_2[0],mul2_out[48][1]);
mul_20x8bit m2_145 (image2[19],filter_2[1],mul2_out[48][2]);
mul_20x8bit m2_146 (image2[20],filter_2[2],mul2_out[48][3]);
mul_20x8bit m2_147 (image2[31],filter_2[3],mul2_out[49][1]);
mul_20x8bit m2_148 (image2[32],filter_2[4],mul2_out[49][2]);
mul_20x8bit m2_149 (image2[33],filter_2[5],mul2_out[49][3]);
mul_20x8bit m2_150 (image2[44],filter_2[6],mul2_out[50][1]);
mul_20x8bit m2_151 (image2[45],filter_2[7],mul2_out[50][2]);
mul_20x8bit m2_152 (image2[46],filter_2[8],mul2_out[50][3]);

adder_24bit ad2_16 (mul2_out[48][1],mul2_out[48][2],mul2_out[48][3],mul2_out[49][1],mul2_out[49][2],mul2_out[49][3],mul2_out[50][1],mul2_out[50][2],mul2_out[50][3],conv2_out[16]);



mul_20x8bit m2_153 (image2[19],filter_2[0],mul2_out[51][1]);
mul_20x8bit m2_154 (image2[20],filter_2[1],mul2_out[51][2]);
mul_20x8bit m2_155 (image2[21],filter_2[2],mul2_out[51][3]);
mul_20x8bit m2_156 (image2[32],filter_2[3],mul2_out[52][1]);
mul_20x8bit m2_157 (image2[33],filter_2[4],mul2_out[52][2]);
mul_20x8bit m2_158 (image2[34],filter_2[5],mul2_out[52][3]);
mul_20x8bit m2_159 (image2[45],filter_2[6],mul2_out[53][1]);
mul_20x8bit m2_160 (image2[46],filter_2[7],mul2_out[53][2]);
mul_20x8bit m2_161 (image2[47],filter_2[8],mul2_out[53][3]);

adder_24bit ad2_17 (mul2_out[51][1],mul2_out[51][2],mul2_out[51][3],mul2_out[52][1],mul2_out[52][2],mul2_out[52][3],mul2_out[53][1],mul2_out[53][2],mul2_out[53][3],conv2_out[17]);



mul_20x8bit m2_162 (image2[20],filter_2[0],mul2_out[54][1]);
mul_20x8bit m2_163 (image2[21],filter_2[1],mul2_out[54][2]);
mul_20x8bit m2_164 (image2[22],filter_2[2],mul2_out[54][3]);
mul_20x8bit m2_165 (image2[33],filter_2[3],mul2_out[55][1]);
mul_20x8bit m2_166 (image2[34],filter_2[4],mul2_out[55][2]);
mul_20x8bit m2_167 (image2[35],filter_2[5],mul2_out[55][3]);
mul_20x8bit m2_168 (image2[46],filter_2[6],mul2_out[56][1]);
mul_20x8bit m2_169 (image2[47],filter_2[7],mul2_out[56][2]);
mul_20x8bit m2_170 (image2[48],filter_2[8],mul2_out[56][3]);

adder_24bit ad2_18 (mul2_out[54][1],mul2_out[54][2],mul2_out[54][3],mul2_out[55][1],mul2_out[55][2],mul2_out[55][3],mul2_out[56][1],mul2_out[56][2],mul2_out[56][3],conv2_out[18]);



mul_20x8bit m2_171 (image2[21],filter_2[0],mul2_out[57][1]);
mul_20x8bit m2_172 (image2[22],filter_2[1],mul2_out[57][2]);
mul_20x8bit m2_173 (image2[23],filter_2[2],mul2_out[57][3]);
mul_20x8bit m2_174 (image2[34],filter_2[3],mul2_out[58][1]);
mul_20x8bit m2_175 (image2[35],filter_2[4],mul2_out[58][2]);
mul_20x8bit m2_176 (image2[36],filter_2[5],mul2_out[58][3]);
mul_20x8bit m2_177 (image2[47],filter_2[6],mul2_out[59][1]);
mul_20x8bit m2_178 (image2[48],filter_2[7],mul2_out[59][2]);
mul_20x8bit m2_179 (image2[49],filter_2[8],mul2_out[59][3]);

adder_24bit ad2_19 (mul2_out[57][1],mul2_out[57][2],mul2_out[57][3],mul2_out[58][1],mul2_out[58][2],mul2_out[58][3],mul2_out[59][1],mul2_out[59][2],mul2_out[59][3],conv2_out[19]);



mul_20x8bit m2_180 (image2[22],filter_2[0],mul2_out[60][1]);
mul_20x8bit m2_181 (image2[23],filter_2[1],mul2_out[60][2]);
mul_20x8bit m2_182 (image2[24],filter_2[2],mul2_out[60][3]);
mul_20x8bit m2_183 (image2[35],filter_2[3],mul2_out[61][1]);
mul_20x8bit m2_184 (image2[36],filter_2[4],mul2_out[61][2]);
mul_20x8bit m2_185 (image2[37],filter_2[5],mul2_out[61][3]);
mul_20x8bit m2_186 (image2[48],filter_2[6],mul2_out[62][1]);
mul_20x8bit m2_187 (image2[49],filter_2[7],mul2_out[62][2]);
mul_20x8bit m2_188 (image2[50],filter_2[8],mul2_out[62][3]);

adder_24bit ad2_20 (mul2_out[60][1],mul2_out[60][2],mul2_out[60][3],mul2_out[61][1],mul2_out[61][2],mul2_out[61][3],mul2_out[62][1],mul2_out[62][2],mul2_out[62][3],conv2_out[20]);



mul_20x8bit m2_189 (image2[23],filter_2[0],mul2_out[63][1]);
mul_20x8bit m2_190 (image2[24],filter_2[1],mul2_out[63][2]);
mul_20x8bit m2_191 (image2[25],filter_2[2],mul2_out[63][3]);
mul_20x8bit m2_192 (image2[36],filter_2[3],mul2_out[64][1]);
mul_20x8bit m2_193 (image2[37],filter_2[4],mul2_out[64][2]);
mul_20x8bit m2_194 (image2[38],filter_2[5],mul2_out[64][3]);
mul_20x8bit m2_195 (image2[49],filter_2[6],mul2_out[65][1]);
mul_20x8bit m2_196 (image2[50],filter_2[7],mul2_out[65][2]);
mul_20x8bit m2_197 (image2[51],filter_2[8],mul2_out[65][3]);

adder_24bit ad2_21 (mul2_out[63][1],mul2_out[63][2],mul2_out[63][3],mul2_out[64][1],mul2_out[64][2],mul2_out[64][3],mul2_out[65][1],mul2_out[65][2],mul2_out[65][3],conv2_out[21]);



mul_20x8bit m2_198 (image2[26],filter_2[0],mul2_out[66][2]);
mul_20x8bit m2_199 (image2[27],filter_2[1],mul2_out[66][3]);
mul_20x8bit m2_200 (image2[28],filter_2[2],mul2_out[66][4]);
mul_20x8bit m2_201 (image2[39],filter_2[3],mul2_out[67][2]);
mul_20x8bit m2_202 (image2[40],filter_2[4],mul2_out[67][3]);
mul_20x8bit m2_203 (image2[41],filter_2[5],mul2_out[67][4]);
mul_20x8bit m2_204 (image2[52],filter_2[6],mul2_out[68][2]);
mul_20x8bit m2_205 (image2[53],filter_2[7],mul2_out[68][3]);
mul_20x8bit m2_206 (image2[54],filter_2[8],mul2_out[68][4]);

adder_24bit ad2_22 (mul2_out[66][2],mul2_out[66][3],mul2_out[66][4],mul2_out[67][2],mul2_out[67][3],mul2_out[67][4],mul2_out[68][2],mul2_out[68][3],mul2_out[68][4],conv2_out[22]);



mul_20x8bit m2_207 (image2[27],filter_2[0],mul2_out[69][2]);
mul_20x8bit m2_208 (image2[28],filter_2[1],mul2_out[69][3]);
mul_20x8bit m2_209 (image2[29],filter_2[2],mul2_out[69][4]);
mul_20x8bit m2_210 (image2[40],filter_2[3],mul2_out[70][2]);
mul_20x8bit m2_211 (image2[41],filter_2[4],mul2_out[70][3]);
mul_20x8bit m2_212 (image2[42],filter_2[5],mul2_out[70][4]);
mul_20x8bit m2_213 (image2[53],filter_2[6],mul2_out[71][2]);
mul_20x8bit m2_214 (image2[54],filter_2[7],mul2_out[71][3]);
mul_20x8bit m2_215 (image2[55],filter_2[8],mul2_out[71][4]);

adder_24bit ad2_23 (mul2_out[69][2],mul2_out[69][3],mul2_out[69][4],mul2_out[70][2],mul2_out[70][3],mul2_out[70][4],mul2_out[71][2],mul2_out[71][3],mul2_out[71][4],conv2_out[23]);



mul_20x8bit m2_216 (image2[28],filter_2[0],mul2_out[72][2]);
mul_20x8bit m2_217 (image2[29],filter_2[1],mul2_out[72][3]);
mul_20x8bit m2_218 (image2[30],filter_2[2],mul2_out[72][4]);
mul_20x8bit m2_219 (image2[41],filter_2[3],mul2_out[73][2]);
mul_20x8bit m2_220 (image2[42],filter_2[4],mul2_out[73][3]);
mul_20x8bit m2_221 (image2[43],filter_2[5],mul2_out[73][4]);
mul_20x8bit m2_222 (image2[54],filter_2[6],mul2_out[74][2]);
mul_20x8bit m2_223 (image2[55],filter_2[7],mul2_out[74][3]);
mul_20x8bit m2_224 (image2[56],filter_2[8],mul2_out[74][4]);

adder_24bit ad2_24 (mul2_out[72][2],mul2_out[72][3],mul2_out[72][4],mul2_out[73][2],mul2_out[73][3],mul2_out[73][4],mul2_out[74][2],mul2_out[74][3],mul2_out[74][4],conv2_out[24]);



mul_20x8bit m2_225 (image2[29],filter_2[0],mul2_out[75][2]);
mul_20x8bit m2_226 (image2[30],filter_2[1],mul2_out[75][3]);
mul_20x8bit m2_227 (image2[31],filter_2[2],mul2_out[75][4]);
mul_20x8bit m2_228 (image2[42],filter_2[3],mul2_out[76][2]);
mul_20x8bit m2_229 (image2[43],filter_2[4],mul2_out[76][3]);
mul_20x8bit m2_230 (image2[44],filter_2[5],mul2_out[76][4]);
mul_20x8bit m2_231 (image2[55],filter_2[6],mul2_out[77][2]);
mul_20x8bit m2_232 (image2[56],filter_2[7],mul2_out[77][3]);
mul_20x8bit m2_233 (image2[57],filter_2[8],mul2_out[77][4]);

adder_24bit ad2_25 (mul2_out[75][2],mul2_out[75][3],mul2_out[75][4],mul2_out[76][2],mul2_out[76][3],mul2_out[76][4],mul2_out[77][2],mul2_out[77][3],mul2_out[77][4],conv2_out[25]);



mul_20x8bit m2_234 (image2[30],filter_2[0],mul2_out[78][2]);
mul_20x8bit m2_235 (image2[31],filter_2[1],mul2_out[78][3]);
mul_20x8bit m2_236 (image2[32],filter_2[2],mul2_out[78][4]);
mul_20x8bit m2_237 (image2[43],filter_2[3],mul2_out[79][2]);
mul_20x8bit m2_238 (image2[44],filter_2[4],mul2_out[79][3]);
mul_20x8bit m2_239 (image2[45],filter_2[5],mul2_out[79][4]);
mul_20x8bit m2_240 (image2[56],filter_2[6],mul2_out[80][2]);
mul_20x8bit m2_241 (image2[57],filter_2[7],mul2_out[80][3]);
mul_20x8bit m2_242 (image2[58],filter_2[8],mul2_out[80][4]);

adder_24bit ad2_26 (mul2_out[78][2],mul2_out[78][3],mul2_out[78][4],mul2_out[79][2],mul2_out[79][3],mul2_out[79][4],mul2_out[80][2],mul2_out[80][3],mul2_out[80][4],conv2_out[26]);



mul_20x8bit m2_243 (image2[31],filter_2[0],mul2_out[81][2]);
mul_20x8bit m2_244 (image2[32],filter_2[1],mul2_out[81][3]);
mul_20x8bit m2_245 (image2[33],filter_2[2],mul2_out[81][4]);
mul_20x8bit m2_246 (image2[44],filter_2[3],mul2_out[82][2]);
mul_20x8bit m2_247 (image2[45],filter_2[4],mul2_out[82][3]);
mul_20x8bit m2_248 (image2[46],filter_2[5],mul2_out[82][4]);
mul_20x8bit m2_249 (image2[57],filter_2[6],mul2_out[83][2]);
mul_20x8bit m2_250 (image2[58],filter_2[7],mul2_out[83][3]);
mul_20x8bit m2_251 (image2[59],filter_2[8],mul2_out[83][4]);

adder_24bit ad2_27 (mul2_out[81][2],mul2_out[81][3],mul2_out[81][4],mul2_out[82][2],mul2_out[82][3],mul2_out[82][4],mul2_out[83][2],mul2_out[83][3],mul2_out[83][4],conv2_out[27]);



mul_20x8bit m2_252 (image2[32],filter_2[0],mul2_out[84][2]);
mul_20x8bit m2_253 (image2[33],filter_2[1],mul2_out[84][3]);
mul_20x8bit m2_254 (image2[34],filter_2[2],mul2_out[84][4]);
mul_20x8bit m2_255 (image2[45],filter_2[3],mul2_out[85][2]);
mul_20x8bit m2_256 (image2[46],filter_2[4],mul2_out[85][3]);
mul_20x8bit m2_257 (image2[47],filter_2[5],mul2_out[85][4]);
mul_20x8bit m2_258 (image2[58],filter_2[6],mul2_out[86][2]);
mul_20x8bit m2_259 (image2[59],filter_2[7],mul2_out[86][3]);
mul_20x8bit m2_260 (image2[60],filter_2[8],mul2_out[86][4]);

adder_24bit ad2_28 (mul2_out[84][2],mul2_out[84][3],mul2_out[84][4],mul2_out[85][2],mul2_out[85][3],mul2_out[85][4],mul2_out[86][2],mul2_out[86][3],mul2_out[86][4],conv2_out[28]);



mul_20x8bit m2_261 (image2[33],filter_2[0],mul2_out[87][2]);
mul_20x8bit m2_262 (image2[34],filter_2[1],mul2_out[87][3]);
mul_20x8bit m2_263 (image2[35],filter_2[2],mul2_out[87][4]);
mul_20x8bit m2_264 (image2[46],filter_2[3],mul2_out[88][2]);
mul_20x8bit m2_265 (image2[47],filter_2[4],mul2_out[88][3]);
mul_20x8bit m2_266 (image2[48],filter_2[5],mul2_out[88][4]);
mul_20x8bit m2_267 (image2[59],filter_2[6],mul2_out[89][2]);
mul_20x8bit m2_268 (image2[60],filter_2[7],mul2_out[89][3]);
mul_20x8bit m2_269 (image2[61],filter_2[8],mul2_out[89][4]);

adder_24bit ad2_29 (mul2_out[87][2],mul2_out[87][3],mul2_out[87][4],mul2_out[88][2],mul2_out[88][3],mul2_out[88][4],mul2_out[89][2],mul2_out[89][3],mul2_out[89][4],conv2_out[29]);



mul_20x8bit m2_270 (image2[34],filter_2[0],mul2_out[90][2]);
mul_20x8bit m2_271 (image2[35],filter_2[1],mul2_out[90][3]);
mul_20x8bit m2_272 (image2[36],filter_2[2],mul2_out[90][4]);
mul_20x8bit m2_273 (image2[47],filter_2[3],mul2_out[91][2]);
mul_20x8bit m2_274 (image2[48],filter_2[4],mul2_out[91][3]);
mul_20x8bit m2_275 (image2[49],filter_2[5],mul2_out[91][4]);
mul_20x8bit m2_276 (image2[60],filter_2[6],mul2_out[92][2]);
mul_20x8bit m2_277 (image2[61],filter_2[7],mul2_out[92][3]);
mul_20x8bit m2_278 (image2[62],filter_2[8],mul2_out[92][4]);

adder_24bit ad2_30 (mul2_out[90][2],mul2_out[90][3],mul2_out[90][4],mul2_out[91][2],mul2_out[91][3],mul2_out[91][4],mul2_out[92][2],mul2_out[92][3],mul2_out[92][4],conv2_out[30]);



mul_20x8bit m2_279 (image2[35],filter_2[0],mul2_out[93][2]);
mul_20x8bit m2_280 (image2[36],filter_2[1],mul2_out[93][3]);
mul_20x8bit m2_281 (image2[37],filter_2[2],mul2_out[93][4]);
mul_20x8bit m2_282 (image2[48],filter_2[3],mul2_out[94][2]);
mul_20x8bit m2_283 (image2[49],filter_2[4],mul2_out[94][3]);
mul_20x8bit m2_284 (image2[50],filter_2[5],mul2_out[94][4]);
mul_20x8bit m2_285 (image2[61],filter_2[6],mul2_out[95][2]);
mul_20x8bit m2_286 (image2[62],filter_2[7],mul2_out[95][3]);
mul_20x8bit m2_287 (image2[63],filter_2[8],mul2_out[95][4]);

adder_24bit ad2_31 (mul2_out[93][2],mul2_out[93][3],mul2_out[93][4],mul2_out[94][2],mul2_out[94][3],mul2_out[94][4],mul2_out[95][2],mul2_out[95][3],mul2_out[95][4],conv2_out[31]);



mul_20x8bit m2_288 (image2[36],filter_2[0],mul2_out[96][2]);
mul_20x8bit m2_289 (image2[37],filter_2[1],mul2_out[96][3]);
mul_20x8bit m2_290 (image2[38],filter_2[2],mul2_out[96][4]);
mul_20x8bit m2_291 (image2[49],filter_2[3],mul2_out[97][2]);
mul_20x8bit m2_292 (image2[50],filter_2[4],mul2_out[97][3]);
mul_20x8bit m2_293 (image2[51],filter_2[5],mul2_out[97][4]);
mul_20x8bit m2_294 (image2[62],filter_2[6],mul2_out[98][2]);
mul_20x8bit m2_295 (image2[63],filter_2[7],mul2_out[98][3]);
mul_20x8bit m2_296 (image2[64],filter_2[8],mul2_out[98][4]);

adder_24bit ad2_32 (mul2_out[96][2],mul2_out[96][3],mul2_out[96][4],mul2_out[97][2],mul2_out[97][3],mul2_out[97][4],mul2_out[98][2],mul2_out[98][3],mul2_out[98][4],conv2_out[32]);



mul_20x8bit m2_297 (image2[39],filter_2[0],mul2_out[99][3]);
mul_20x8bit m2_298 (image2[40],filter_2[1],mul2_out[99][4]);
mul_20x8bit m2_299 (image2[41],filter_2[2],mul2_out[99][5]);
mul_20x8bit m2_300 (image2[52],filter_2[3],mul2_out[100][3]);
mul_20x8bit m2_301 (image2[53],filter_2[4],mul2_out[100][4]);
mul_20x8bit m2_302 (image2[54],filter_2[5],mul2_out[100][5]);
mul_20x8bit m2_303 (image2[65],filter_2[6],mul2_out[101][3]);
mul_20x8bit m2_304 (image2[66],filter_2[7],mul2_out[101][4]);
mul_20x8bit m2_305 (image2[67],filter_2[8],mul2_out[101][5]);

adder_24bit ad2_33 (mul2_out[99][3],mul2_out[99][4],mul2_out[99][5],mul2_out[100][3],mul2_out[100][4],mul2_out[100][5],mul2_out[101][3],mul2_out[101][4],mul2_out[101][5],conv2_out[33]);



mul_20x8bit m2_306 (image2[40],filter_2[0],mul2_out[102][3]);
mul_20x8bit m2_307 (image2[41],filter_2[1],mul2_out[102][4]);
mul_20x8bit m2_308 (image2[42],filter_2[2],mul2_out[102][5]);
mul_20x8bit m2_309 (image2[53],filter_2[3],mul2_out[103][3]);
mul_20x8bit m2_310 (image2[54],filter_2[4],mul2_out[103][4]);
mul_20x8bit m2_311 (image2[55],filter_2[5],mul2_out[103][5]);
mul_20x8bit m2_312 (image2[66],filter_2[6],mul2_out[104][3]);
mul_20x8bit m2_313 (image2[67],filter_2[7],mul2_out[104][4]);
mul_20x8bit m2_314 (image2[68],filter_2[8],mul2_out[104][5]);

adder_24bit ad2_34 (mul2_out[102][3],mul2_out[102][4],mul2_out[102][5],mul2_out[103][3],mul2_out[103][4],mul2_out[103][5],mul2_out[104][3],mul2_out[104][4],mul2_out[104][5],conv2_out[34]);



mul_20x8bit m2_315 (image2[41],filter_2[0],mul2_out[105][3]);
mul_20x8bit m2_316 (image2[42],filter_2[1],mul2_out[105][4]);
mul_20x8bit m2_317 (image2[43],filter_2[2],mul2_out[105][5]);
mul_20x8bit m2_318 (image2[54],filter_2[3],mul2_out[106][3]);
mul_20x8bit m2_319 (image2[55],filter_2[4],mul2_out[106][4]);
mul_20x8bit m2_320 (image2[56],filter_2[5],mul2_out[106][5]);
mul_20x8bit m2_321 (image2[67],filter_2[6],mul2_out[107][3]);
mul_20x8bit m2_322 (image2[68],filter_2[7],mul2_out[107][4]);
mul_20x8bit m2_323 (image2[69],filter_2[8],mul2_out[107][5]);

adder_24bit ad2_35 (mul2_out[105][3],mul2_out[105][4],mul2_out[105][5],mul2_out[106][3],mul2_out[106][4],mul2_out[106][5],mul2_out[107][3],mul2_out[107][4],mul2_out[107][5],conv2_out[35]);



mul_20x8bit m2_324 (image2[42],filter_2[0],mul2_out[108][3]);
mul_20x8bit m2_325 (image2[43],filter_2[1],mul2_out[108][4]);
mul_20x8bit m2_326 (image2[44],filter_2[2],mul2_out[108][5]);
mul_20x8bit m2_327 (image2[55],filter_2[3],mul2_out[109][3]);
mul_20x8bit m2_328 (image2[56],filter_2[4],mul2_out[109][4]);
mul_20x8bit m2_329 (image2[57],filter_2[5],mul2_out[109][5]);
mul_20x8bit m2_330 (image2[68],filter_2[6],mul2_out[110][3]);
mul_20x8bit m2_331 (image2[69],filter_2[7],mul2_out[110][4]);
mul_20x8bit m2_332 (image2[70],filter_2[8],mul2_out[110][5]);

adder_24bit ad2_36 (mul2_out[108][3],mul2_out[108][4],mul2_out[108][5],mul2_out[109][3],mul2_out[109][4],mul2_out[109][5],mul2_out[110][3],mul2_out[110][4],mul2_out[110][5],conv2_out[36]);



mul_20x8bit m2_333 (image2[43],filter_2[0],mul2_out[111][3]);
mul_20x8bit m2_334 (image2[44],filter_2[1],mul2_out[111][4]);
mul_20x8bit m2_335 (image2[45],filter_2[2],mul2_out[111][5]);
mul_20x8bit m2_336 (image2[56],filter_2[3],mul2_out[112][3]);
mul_20x8bit m2_337 (image2[57],filter_2[4],mul2_out[112][4]);
mul_20x8bit m2_338 (image2[58],filter_2[5],mul2_out[112][5]);
mul_20x8bit m2_339 (image2[69],filter_2[6],mul2_out[113][3]);
mul_20x8bit m2_340 (image2[70],filter_2[7],mul2_out[113][4]);
mul_20x8bit m2_341 (image2[71],filter_2[8],mul2_out[113][5]);

adder_24bit ad2_37 (mul2_out[111][3],mul2_out[111][4],mul2_out[111][5],mul2_out[112][3],mul2_out[112][4],mul2_out[112][5],mul2_out[113][3],mul2_out[113][4],mul2_out[113][5],conv2_out[37]);



mul_20x8bit m2_342 (image2[44],filter_2[0],mul2_out[114][3]);
mul_20x8bit m2_343 (image2[45],filter_2[1],mul2_out[114][4]);
mul_20x8bit m2_344 (image2[46],filter_2[2],mul2_out[114][5]);
mul_20x8bit m2_345 (image2[57],filter_2[3],mul2_out[115][3]);
mul_20x8bit m2_346 (image2[58],filter_2[4],mul2_out[115][4]);
mul_20x8bit m2_347 (image2[59],filter_2[5],mul2_out[115][5]);
mul_20x8bit m2_348 (image2[70],filter_2[6],mul2_out[116][3]);
mul_20x8bit m2_349 (image2[71],filter_2[7],mul2_out[116][4]);
mul_20x8bit m2_350 (image2[72],filter_2[8],mul2_out[116][5]);

adder_24bit ad2_38 (mul2_out[114][3],mul2_out[114][4],mul2_out[114][5],mul2_out[115][3],mul2_out[115][4],mul2_out[115][5],mul2_out[116][3],mul2_out[116][4],mul2_out[116][5],conv2_out[38]);



mul_20x8bit m2_351 (image2[45],filter_2[0],mul2_out[117][3]);
mul_20x8bit m2_352 (image2[46],filter_2[1],mul2_out[117][4]);
mul_20x8bit m2_353 (image2[47],filter_2[2],mul2_out[117][5]);
mul_20x8bit m2_354 (image2[58],filter_2[3],mul2_out[118][3]);
mul_20x8bit m2_355 (image2[59],filter_2[4],mul2_out[118][4]);
mul_20x8bit m2_356 (image2[60],filter_2[5],mul2_out[118][5]);
mul_20x8bit m2_357 (image2[71],filter_2[6],mul2_out[119][3]);
mul_20x8bit m2_358 (image2[72],filter_2[7],mul2_out[119][4]);
mul_20x8bit m2_359 (image2[73],filter_2[8],mul2_out[119][5]);

adder_24bit ad2_39 (mul2_out[117][3],mul2_out[117][4],mul2_out[117][5],mul2_out[118][3],mul2_out[118][4],mul2_out[118][5],mul2_out[119][3],mul2_out[119][4],mul2_out[119][5],conv2_out[39]);



mul_20x8bit m2_360 (image2[46],filter_2[0],mul2_out[120][3]);
mul_20x8bit m2_361 (image2[47],filter_2[1],mul2_out[120][4]);
mul_20x8bit m2_362 (image2[48],filter_2[2],mul2_out[120][5]);
mul_20x8bit m2_363 (image2[59],filter_2[3],mul2_out[121][3]);
mul_20x8bit m2_364 (image2[60],filter_2[4],mul2_out[121][4]);
mul_20x8bit m2_365 (image2[61],filter_2[5],mul2_out[121][5]);
mul_20x8bit m2_366 (image2[72],filter_2[6],mul2_out[122][3]);
mul_20x8bit m2_367 (image2[73],filter_2[7],mul2_out[122][4]);
mul_20x8bit m2_368 (image2[74],filter_2[8],mul2_out[122][5]);

adder_24bit ad2_40 (mul2_out[120][3],mul2_out[120][4],mul2_out[120][5],mul2_out[121][3],mul2_out[121][4],mul2_out[121][5],mul2_out[122][3],mul2_out[122][4],mul2_out[122][5],conv2_out[40]);



mul_20x8bit m2_369 (image2[47],filter_2[0],mul2_out[123][3]);
mul_20x8bit m2_370 (image2[48],filter_2[1],mul2_out[123][4]);
mul_20x8bit m2_371 (image2[49],filter_2[2],mul2_out[123][5]);
mul_20x8bit m2_372 (image2[60],filter_2[3],mul2_out[124][3]);
mul_20x8bit m2_373 (image2[61],filter_2[4],mul2_out[124][4]);
mul_20x8bit m2_374 (image2[62],filter_2[5],mul2_out[124][5]);
mul_20x8bit m2_375 (image2[73],filter_2[6],mul2_out[125][3]);
mul_20x8bit m2_376 (image2[74],filter_2[7],mul2_out[125][4]);
mul_20x8bit m2_377 (image2[75],filter_2[8],mul2_out[125][5]);

adder_24bit ad2_41 (mul2_out[123][3],mul2_out[123][4],mul2_out[123][5],mul2_out[124][3],mul2_out[124][4],mul2_out[124][5],mul2_out[125][3],mul2_out[125][4],mul2_out[125][5],conv2_out[41]);



mul_20x8bit m2_378 (image2[48],filter_2[0],mul2_out[126][3]);
mul_20x8bit m2_379 (image2[49],filter_2[1],mul2_out[126][4]);
mul_20x8bit m2_380 (image2[50],filter_2[2],mul2_out[126][5]);
mul_20x8bit m2_381 (image2[61],filter_2[3],mul2_out[127][3]);
mul_20x8bit m2_382 (image2[62],filter_2[4],mul2_out[127][4]);
mul_20x8bit m2_383 (image2[63],filter_2[5],mul2_out[127][5]);
mul_20x8bit m2_384 (image2[74],filter_2[6],mul2_out[128][3]);
mul_20x8bit m2_385 (image2[75],filter_2[7],mul2_out[128][4]);
mul_20x8bit m2_386 (image2[76],filter_2[8],mul2_out[128][5]);

adder_24bit ad2_42 (mul2_out[126][3],mul2_out[126][4],mul2_out[126][5],mul2_out[127][3],mul2_out[127][4],mul2_out[127][5],mul2_out[128][3],mul2_out[128][4],mul2_out[128][5],conv2_out[42]);



mul_20x8bit m2_387 (image2[49],filter_2[0],mul2_out[129][3]);
mul_20x8bit m2_388 (image2[50],filter_2[1],mul2_out[129][4]);
mul_20x8bit m2_389 (image2[51],filter_2[2],mul2_out[129][5]);
mul_20x8bit m2_390 (image2[62],filter_2[3],mul2_out[130][3]);
mul_20x8bit m2_391 (image2[63],filter_2[4],mul2_out[130][4]);
mul_20x8bit m2_392 (image2[64],filter_2[5],mul2_out[130][5]);
mul_20x8bit m2_393 (image2[75],filter_2[6],mul2_out[131][3]);
mul_20x8bit m2_394 (image2[76],filter_2[7],mul2_out[131][4]);
mul_20x8bit m2_395 (image2[77],filter_2[8],mul2_out[131][5]);

adder_24bit ad2_43 (mul2_out[129][3],mul2_out[129][4],mul2_out[129][5],mul2_out[130][3],mul2_out[130][4],mul2_out[130][5],mul2_out[131][3],mul2_out[131][4],mul2_out[131][5],conv2_out[43]);



mul_20x8bit m2_396 (image2[52],filter_2[0],mul2_out[132][4]);
mul_20x8bit m2_397 (image2[53],filter_2[1],mul2_out[132][5]);
mul_20x8bit m2_398 (image2[54],filter_2[2],mul2_out[132][6]);
mul_20x8bit m2_399 (image2[65],filter_2[3],mul2_out[133][4]);
mul_20x8bit m2_400 (image2[66],filter_2[4],mul2_out[133][5]);
mul_20x8bit m2_401 (image2[67],filter_2[5],mul2_out[133][6]);
mul_20x8bit m2_402 (image2[78],filter_2[6],mul2_out[134][4]);
mul_20x8bit m2_403 (image2[79],filter_2[7],mul2_out[134][5]);
mul_20x8bit m2_404 (image2[80],filter_2[8],mul2_out[134][6]);

adder_24bit ad2_44 (mul2_out[132][4],mul2_out[132][5],mul2_out[132][6],mul2_out[133][4],mul2_out[133][5],mul2_out[133][6],mul2_out[134][4],mul2_out[134][5],mul2_out[134][6],conv2_out[44]);



mul_20x8bit m2_405 (image2[53],filter_2[0],mul2_out[135][4]);
mul_20x8bit m2_406 (image2[54],filter_2[1],mul2_out[135][5]);
mul_20x8bit m2_407 (image2[55],filter_2[2],mul2_out[135][6]);
mul_20x8bit m2_408 (image2[66],filter_2[3],mul2_out[136][4]);
mul_20x8bit m2_409 (image2[67],filter_2[4],mul2_out[136][5]);
mul_20x8bit m2_410 (image2[68],filter_2[5],mul2_out[136][6]);
mul_20x8bit m2_411 (image2[79],filter_2[6],mul2_out[137][4]);
mul_20x8bit m2_412 (image2[80],filter_2[7],mul2_out[137][5]);
mul_20x8bit m2_413 (image2[81],filter_2[8],mul2_out[137][6]);

adder_24bit ad2_45 (mul2_out[135][4],mul2_out[135][5],mul2_out[135][6],mul2_out[136][4],mul2_out[136][5],mul2_out[136][6],mul2_out[137][4],mul2_out[137][5],mul2_out[137][6],conv2_out[45]);



mul_20x8bit m2_414 (image2[54],filter_2[0],mul2_out[138][4]);
mul_20x8bit m2_415 (image2[55],filter_2[1],mul2_out[138][5]);
mul_20x8bit m2_416 (image2[56],filter_2[2],mul2_out[138][6]);
mul_20x8bit m2_417 (image2[67],filter_2[3],mul2_out[139][4]);
mul_20x8bit m2_418 (image2[68],filter_2[4],mul2_out[139][5]);
mul_20x8bit m2_419 (image2[69],filter_2[5],mul2_out[139][6]);
mul_20x8bit m2_420 (image2[80],filter_2[6],mul2_out[140][4]);
mul_20x8bit m2_421 (image2[81],filter_2[7],mul2_out[140][5]);
mul_20x8bit m2_422 (image2[82],filter_2[8],mul2_out[140][6]);

adder_24bit ad2_46 (mul2_out[138][4],mul2_out[138][5],mul2_out[138][6],mul2_out[139][4],mul2_out[139][5],mul2_out[139][6],mul2_out[140][4],mul2_out[140][5],mul2_out[140][6],conv2_out[46]);



mul_20x8bit m2_423 (image2[55],filter_2[0],mul2_out[141][4]);
mul_20x8bit m2_424 (image2[56],filter_2[1],mul2_out[141][5]);
mul_20x8bit m2_425 (image2[57],filter_2[2],mul2_out[141][6]);
mul_20x8bit m2_426 (image2[68],filter_2[3],mul2_out[142][4]);
mul_20x8bit m2_427 (image2[69],filter_2[4],mul2_out[142][5]);
mul_20x8bit m2_428 (image2[70],filter_2[5],mul2_out[142][6]);
mul_20x8bit m2_429 (image2[81],filter_2[6],mul2_out[143][4]);
mul_20x8bit m2_430 (image2[82],filter_2[7],mul2_out[143][5]);
mul_20x8bit m2_431 (image2[83],filter_2[8],mul2_out[143][6]);

adder_24bit ad2_47 (mul2_out[141][4],mul2_out[141][5],mul2_out[141][6],mul2_out[142][4],mul2_out[142][5],mul2_out[142][6],mul2_out[143][4],mul2_out[143][5],mul2_out[143][6],conv2_out[47]);



mul_20x8bit m2_432 (image2[56],filter_2[0],mul2_out[144][4]);
mul_20x8bit m2_433 (image2[57],filter_2[1],mul2_out[144][5]);
mul_20x8bit m2_434 (image2[58],filter_2[2],mul2_out[144][6]);
mul_20x8bit m2_435 (image2[69],filter_2[3],mul2_out[145][4]);
mul_20x8bit m2_436 (image2[70],filter_2[4],mul2_out[145][5]);
mul_20x8bit m2_437 (image2[71],filter_2[5],mul2_out[145][6]);
mul_20x8bit m2_438 (image2[82],filter_2[6],mul2_out[146][4]);
mul_20x8bit m2_439 (image2[83],filter_2[7],mul2_out[146][5]);
mul_20x8bit m2_440 (image2[84],filter_2[8],mul2_out[146][6]);

adder_24bit ad2_48 (mul2_out[144][4],mul2_out[144][5],mul2_out[144][6],mul2_out[145][4],mul2_out[145][5],mul2_out[145][6],mul2_out[146][4],mul2_out[146][5],mul2_out[146][6],conv2_out[48]);



mul_20x8bit m2_441 (image2[57],filter_2[0],mul2_out[147][4]);
mul_20x8bit m2_442 (image2[58],filter_2[1],mul2_out[147][5]);
mul_20x8bit m2_443 (image2[59],filter_2[2],mul2_out[147][6]);
mul_20x8bit m2_444 (image2[70],filter_2[3],mul2_out[148][4]);
mul_20x8bit m2_445 (image2[71],filter_2[4],mul2_out[148][5]);
mul_20x8bit m2_446 (image2[72],filter_2[5],mul2_out[148][6]);
mul_20x8bit m2_447 (image2[83],filter_2[6],mul2_out[149][4]);
mul_20x8bit m2_448 (image2[84],filter_2[7],mul2_out[149][5]);
mul_20x8bit m2_449 (image2[85],filter_2[8],mul2_out[149][6]);

adder_24bit ad2_49 (mul2_out[147][4],mul2_out[147][5],mul2_out[147][6],mul2_out[148][4],mul2_out[148][5],mul2_out[148][6],mul2_out[149][4],mul2_out[149][5],mul2_out[149][6],conv2_out[49]);



mul_20x8bit m2_450 (image2[58],filter_2[0],mul2_out[150][4]);
mul_20x8bit m2_451 (image2[59],filter_2[1],mul2_out[150][5]);
mul_20x8bit m2_452 (image2[60],filter_2[2],mul2_out[150][6]);
mul_20x8bit m2_453 (image2[71],filter_2[3],mul2_out[151][4]);
mul_20x8bit m2_454 (image2[72],filter_2[4],mul2_out[151][5]);
mul_20x8bit m2_455 (image2[73],filter_2[5],mul2_out[151][6]);
mul_20x8bit m2_456 (image2[84],filter_2[6],mul2_out[152][4]);
mul_20x8bit m2_457 (image2[85],filter_2[7],mul2_out[152][5]);
mul_20x8bit m2_458 (image2[86],filter_2[8],mul2_out[152][6]);

adder_24bit ad2_50 (mul2_out[150][4],mul2_out[150][5],mul2_out[150][6],mul2_out[151][4],mul2_out[151][5],mul2_out[151][6],mul2_out[152][4],mul2_out[152][5],mul2_out[152][6],conv2_out[50]);



mul_20x8bit m2_459 (image2[59],filter_2[0],mul2_out[153][4]);
mul_20x8bit m2_460 (image2[60],filter_2[1],mul2_out[153][5]);
mul_20x8bit m2_461 (image2[61],filter_2[2],mul2_out[153][6]);
mul_20x8bit m2_462 (image2[72],filter_2[3],mul2_out[154][4]);
mul_20x8bit m2_463 (image2[73],filter_2[4],mul2_out[154][5]);
mul_20x8bit m2_464 (image2[74],filter_2[5],mul2_out[154][6]);
mul_20x8bit m2_465 (image2[85],filter_2[6],mul2_out[155][4]);
mul_20x8bit m2_466 (image2[86],filter_2[7],mul2_out[155][5]);
mul_20x8bit m2_467 (image2[87],filter_2[8],mul2_out[155][6]);

adder_24bit ad2_51 (mul2_out[153][4],mul2_out[153][5],mul2_out[153][6],mul2_out[154][4],mul2_out[154][5],mul2_out[154][6],mul2_out[155][4],mul2_out[155][5],mul2_out[155][6],conv2_out[51]);



mul_20x8bit m2_468 (image2[60],filter_2[0],mul2_out[156][4]);
mul_20x8bit m2_469 (image2[61],filter_2[1],mul2_out[156][5]);
mul_20x8bit m2_470 (image2[62],filter_2[2],mul2_out[156][6]);
mul_20x8bit m2_471 (image2[73],filter_2[3],mul2_out[157][4]);
mul_20x8bit m2_472 (image2[74],filter_2[4],mul2_out[157][5]);
mul_20x8bit m2_473 (image2[75],filter_2[5],mul2_out[157][6]);
mul_20x8bit m2_474 (image2[86],filter_2[6],mul2_out[158][4]);
mul_20x8bit m2_475 (image2[87],filter_2[7],mul2_out[158][5]);
mul_20x8bit m2_476 (image2[88],filter_2[8],mul2_out[158][6]);

adder_24bit ad2_52 (mul2_out[156][4],mul2_out[156][5],mul2_out[156][6],mul2_out[157][4],mul2_out[157][5],mul2_out[157][6],mul2_out[158][4],mul2_out[158][5],mul2_out[158][6],conv2_out[52]);



mul_20x8bit m2_477 (image2[61],filter_2[0],mul2_out[159][4]);
mul_20x8bit m2_478 (image2[62],filter_2[1],mul2_out[159][5]);
mul_20x8bit m2_479 (image2[63],filter_2[2],mul2_out[159][6]);
mul_20x8bit m2_480 (image2[74],filter_2[3],mul2_out[160][4]);
mul_20x8bit m2_481 (image2[75],filter_2[4],mul2_out[160][5]);
mul_20x8bit m2_482 (image2[76],filter_2[5],mul2_out[160][6]);
mul_20x8bit m2_483 (image2[87],filter_2[6],mul2_out[161][4]);
mul_20x8bit m2_484 (image2[88],filter_2[7],mul2_out[161][5]);
mul_20x8bit m2_485 (image2[89],filter_2[8],mul2_out[161][6]);

adder_24bit ad2_53 (mul2_out[159][4],mul2_out[159][5],mul2_out[159][6],mul2_out[160][4],mul2_out[160][5],mul2_out[160][6],mul2_out[161][4],mul2_out[161][5],mul2_out[161][6],conv2_out[53]);



mul_20x8bit m2_486 (image2[62],filter_2[0],mul2_out[162][4]);
mul_20x8bit m2_487 (image2[63],filter_2[1],mul2_out[162][5]);
mul_20x8bit m2_488 (image2[64],filter_2[2],mul2_out[162][6]);
mul_20x8bit m2_489 (image2[75],filter_2[3],mul2_out[163][4]);
mul_20x8bit m2_490 (image2[76],filter_2[4],mul2_out[163][5]);
mul_20x8bit m2_491 (image2[77],filter_2[5],mul2_out[163][6]);
mul_20x8bit m2_492 (image2[88],filter_2[6],mul2_out[164][4]);
mul_20x8bit m2_493 (image2[89],filter_2[7],mul2_out[164][5]);
mul_20x8bit m2_494 (image2[90],filter_2[8],mul2_out[164][6]);

adder_24bit ad2_54 (mul2_out[162][4],mul2_out[162][5],mul2_out[162][6],mul2_out[163][4],mul2_out[163][5],mul2_out[163][6],mul2_out[164][4],mul2_out[164][5],mul2_out[164][6],conv2_out[54]);



mul_20x8bit m2_495 (image2[65],filter_2[0],mul2_out[165][5]);
mul_20x8bit m2_496 (image2[66],filter_2[1],mul2_out[165][6]);
mul_20x8bit m2_497 (image2[67],filter_2[2],mul2_out[165][7]);
mul_20x8bit m2_498 (image2[78],filter_2[3],mul2_out[166][5]);
mul_20x8bit m2_499 (image2[79],filter_2[4],mul2_out[166][6]);
mul_20x8bit m2_500 (image2[80],filter_2[5],mul2_out[166][7]);
mul_20x8bit m2_501 (image2[91],filter_2[6],mul2_out[167][5]);
mul_20x8bit m2_502 (image2[92],filter_2[7],mul2_out[167][6]);
mul_20x8bit m2_503 (image2[93],filter_2[8],mul2_out[167][7]);

adder_24bit ad2_55 (mul2_out[165][5],mul2_out[165][6],mul2_out[165][7],mul2_out[166][5],mul2_out[166][6],mul2_out[166][7],mul2_out[167][5],mul2_out[167][6],mul2_out[167][7],conv2_out[55]);



mul_20x8bit m2_504 (image2[66],filter_2[0],mul2_out[168][5]);
mul_20x8bit m2_505 (image2[67],filter_2[1],mul2_out[168][6]);
mul_20x8bit m2_506 (image2[68],filter_2[2],mul2_out[168][7]);
mul_20x8bit m2_507 (image2[79],filter_2[3],mul2_out[169][5]);
mul_20x8bit m2_508 (image2[80],filter_2[4],mul2_out[169][6]);
mul_20x8bit m2_509 (image2[81],filter_2[5],mul2_out[169][7]);
mul_20x8bit m2_510 (image2[92],filter_2[6],mul2_out[170][5]);
mul_20x8bit m2_511 (image2[93],filter_2[7],mul2_out[170][6]);
mul_20x8bit m2_512 (image2[94],filter_2[8],mul2_out[170][7]);

adder_24bit ad2_56 (mul2_out[168][5],mul2_out[168][6],mul2_out[168][7],mul2_out[169][5],mul2_out[169][6],mul2_out[169][7],mul2_out[170][5],mul2_out[170][6],mul2_out[170][7],conv2_out[56]);



mul_20x8bit m2_513 (image2[67],filter_2[0],mul2_out[171][5]);
mul_20x8bit m2_514 (image2[68],filter_2[1],mul2_out[171][6]);
mul_20x8bit m2_515 (image2[69],filter_2[2],mul2_out[171][7]);
mul_20x8bit m2_516 (image2[80],filter_2[3],mul2_out[172][5]);
mul_20x8bit m2_517 (image2[81],filter_2[4],mul2_out[172][6]);
mul_20x8bit m2_518 (image2[82],filter_2[5],mul2_out[172][7]);
mul_20x8bit m2_519 (image2[93],filter_2[6],mul2_out[173][5]);
mul_20x8bit m2_520 (image2[94],filter_2[7],mul2_out[173][6]);
mul_20x8bit m2_521 (image2[95],filter_2[8],mul2_out[173][7]);

adder_24bit ad2_57 (mul2_out[171][5],mul2_out[171][6],mul2_out[171][7],mul2_out[172][5],mul2_out[172][6],mul2_out[172][7],mul2_out[173][5],mul2_out[173][6],mul2_out[173][7],conv2_out[57]);



mul_20x8bit m2_522 (image2[68],filter_2[0],mul2_out[174][5]);
mul_20x8bit m2_523 (image2[69],filter_2[1],mul2_out[174][6]);
mul_20x8bit m2_524 (image2[70],filter_2[2],mul2_out[174][7]);
mul_20x8bit m2_525 (image2[81],filter_2[3],mul2_out[175][5]);
mul_20x8bit m2_526 (image2[82],filter_2[4],mul2_out[175][6]);
mul_20x8bit m2_527 (image2[83],filter_2[5],mul2_out[175][7]);
mul_20x8bit m2_528 (image2[94],filter_2[6],mul2_out[176][5]);
mul_20x8bit m2_529 (image2[95],filter_2[7],mul2_out[176][6]);
mul_20x8bit m2_530 (image2[96],filter_2[8],mul2_out[176][7]);

adder_24bit ad2_58 (mul2_out[174][5],mul2_out[174][6],mul2_out[174][7],mul2_out[175][5],mul2_out[175][6],mul2_out[175][7],mul2_out[176][5],mul2_out[176][6],mul2_out[176][7],conv2_out[58]);



mul_20x8bit m2_531 (image2[69],filter_2[0],mul2_out[177][5]);
mul_20x8bit m2_532 (image2[70],filter_2[1],mul2_out[177][6]);
mul_20x8bit m2_533 (image2[71],filter_2[2],mul2_out[177][7]);
mul_20x8bit m2_534 (image2[82],filter_2[3],mul2_out[178][5]);
mul_20x8bit m2_535 (image2[83],filter_2[4],mul2_out[178][6]);
mul_20x8bit m2_536 (image2[84],filter_2[5],mul2_out[178][7]);
mul_20x8bit m2_537 (image2[95],filter_2[6],mul2_out[179][5]);
mul_20x8bit m2_538 (image2[96],filter_2[7],mul2_out[179][6]);
mul_20x8bit m2_539 (image2[97],filter_2[8],mul2_out[179][7]);

adder_24bit ad2_59 (mul2_out[177][5],mul2_out[177][6],mul2_out[177][7],mul2_out[178][5],mul2_out[178][6],mul2_out[178][7],mul2_out[179][5],mul2_out[179][6],mul2_out[179][7],conv2_out[59]);



mul_20x8bit m2_540 (image2[70],filter_2[0],mul2_out[180][5]);
mul_20x8bit m2_541 (image2[71],filter_2[1],mul2_out[180][6]);
mul_20x8bit m2_542 (image2[72],filter_2[2],mul2_out[180][7]);
mul_20x8bit m2_543 (image2[83],filter_2[3],mul2_out[181][5]);
mul_20x8bit m2_544 (image2[84],filter_2[4],mul2_out[181][6]);
mul_20x8bit m2_545 (image2[85],filter_2[5],mul2_out[181][7]);
mul_20x8bit m2_546 (image2[96],filter_2[6],mul2_out[182][5]);
mul_20x8bit m2_547 (image2[97],filter_2[7],mul2_out[182][6]);
mul_20x8bit m2_548 (image2[98],filter_2[8],mul2_out[182][7]);

adder_24bit ad2_60 (mul2_out[180][5],mul2_out[180][6],mul2_out[180][7],mul2_out[181][5],mul2_out[181][6],mul2_out[181][7],mul2_out[182][5],mul2_out[182][6],mul2_out[182][7],conv2_out[60]);



mul_20x8bit m2_549 (image2[71],filter_2[0],mul2_out[183][5]);
mul_20x8bit m2_550 (image2[72],filter_2[1],mul2_out[183][6]);
mul_20x8bit m2_551 (image2[73],filter_2[2],mul2_out[183][7]);
mul_20x8bit m2_552 (image2[84],filter_2[3],mul2_out[184][5]);
mul_20x8bit m2_553 (image2[85],filter_2[4],mul2_out[184][6]);
mul_20x8bit m2_554 (image2[86],filter_2[5],mul2_out[184][7]);
mul_20x8bit m2_555 (image2[97],filter_2[6],mul2_out[185][5]);
mul_20x8bit m2_556 (image2[98],filter_2[7],mul2_out[185][6]);
mul_20x8bit m2_557 (image2[99],filter_2[8],mul2_out[185][7]);

adder_24bit ad2_61 (mul2_out[183][5],mul2_out[183][6],mul2_out[183][7],mul2_out[184][5],mul2_out[184][6],mul2_out[184][7],mul2_out[185][5],mul2_out[185][6],mul2_out[185][7],conv2_out[61]);



mul_20x8bit m2_558 (image2[72],filter_2[0],mul2_out[186][5]);
mul_20x8bit m2_559 (image2[73],filter_2[1],mul2_out[186][6]);
mul_20x8bit m2_560 (image2[74],filter_2[2],mul2_out[186][7]);
mul_20x8bit m2_561 (image2[85],filter_2[3],mul2_out[187][5]);
mul_20x8bit m2_562 (image2[86],filter_2[4],mul2_out[187][6]);
mul_20x8bit m2_563 (image2[87],filter_2[5],mul2_out[187][7]);
mul_20x8bit m2_564 (image2[98],filter_2[6],mul2_out[188][5]);
mul_20x8bit m2_565 (image2[99],filter_2[7],mul2_out[188][6]);
mul_20x8bit m2_566 (image2[100],filter_2[8],mul2_out[188][7]);

adder_24bit ad2_62 (mul2_out[186][5],mul2_out[186][6],mul2_out[186][7],mul2_out[187][5],mul2_out[187][6],mul2_out[187][7],mul2_out[188][5],mul2_out[188][6],mul2_out[188][7],conv2_out[62]);



mul_20x8bit m2_567 (image2[73],filter_2[0],mul2_out[189][5]);
mul_20x8bit m2_568 (image2[74],filter_2[1],mul2_out[189][6]);
mul_20x8bit m2_569 (image2[75],filter_2[2],mul2_out[189][7]);
mul_20x8bit m2_570 (image2[86],filter_2[3],mul2_out[190][5]);
mul_20x8bit m2_571 (image2[87],filter_2[4],mul2_out[190][6]);
mul_20x8bit m2_572 (image2[88],filter_2[5],mul2_out[190][7]);
mul_20x8bit m2_573 (image2[99],filter_2[6],mul2_out[191][5]);
mul_20x8bit m2_574 (image2[100],filter_2[7],mul2_out[191][6]);
mul_20x8bit m2_575 (image2[101],filter_2[8],mul2_out[191][7]);

adder_24bit ad2_63 (mul2_out[189][5],mul2_out[189][6],mul2_out[189][7],mul2_out[190][5],mul2_out[190][6],mul2_out[190][7],mul2_out[191][5],mul2_out[191][6],mul2_out[191][7],conv2_out[63]);



mul_20x8bit m2_576 (image2[74],filter_2[0],mul2_out[192][5]);
mul_20x8bit m2_577 (image2[75],filter_2[1],mul2_out[192][6]);
mul_20x8bit m2_578 (image2[76],filter_2[2],mul2_out[192][7]);
mul_20x8bit m2_579 (image2[87],filter_2[3],mul2_out[193][5]);
mul_20x8bit m2_580 (image2[88],filter_2[4],mul2_out[193][6]);
mul_20x8bit m2_581 (image2[89],filter_2[5],mul2_out[193][7]);
mul_20x8bit m2_582 (image2[100],filter_2[6],mul2_out[194][5]);
mul_20x8bit m2_583 (image2[101],filter_2[7],mul2_out[194][6]);
mul_20x8bit m2_584 (image2[102],filter_2[8],mul2_out[194][7]);

adder_24bit ad2_64 (mul2_out[192][5],mul2_out[192][6],mul2_out[192][7],mul2_out[193][5],mul2_out[193][6],mul2_out[193][7],mul2_out[194][5],mul2_out[194][6],mul2_out[194][7],conv2_out[64]);



mul_20x8bit m2_585 (image2[75],filter_2[0],mul2_out[195][5]);
mul_20x8bit m2_586 (image2[76],filter_2[1],mul2_out[195][6]);
mul_20x8bit m2_587 (image2[77],filter_2[2],mul2_out[195][7]);
mul_20x8bit m2_588 (image2[88],filter_2[3],mul2_out[196][5]);
mul_20x8bit m2_589 (image2[89],filter_2[4],mul2_out[196][6]);
mul_20x8bit m2_590 (image2[90],filter_2[5],mul2_out[196][7]);
mul_20x8bit m2_591 (image2[101],filter_2[6],mul2_out[197][5]);
mul_20x8bit m2_592 (image2[102],filter_2[7],mul2_out[197][6]);
mul_20x8bit m2_593 (image2[103],filter_2[8],mul2_out[197][7]);

adder_24bit ad2_65 (mul2_out[195][5],mul2_out[195][6],mul2_out[195][7],mul2_out[196][5],mul2_out[196][6],mul2_out[196][7],mul2_out[197][5],mul2_out[197][6],mul2_out[197][7],conv2_out[65]);



mul_20x8bit m2_594 (image2[78],filter_2[0],mul2_out[198][6]);
mul_20x8bit m2_595 (image2[79],filter_2[1],mul2_out[198][7]);
mul_20x8bit m2_596 (image2[80],filter_2[2],mul2_out[198][8]);
mul_20x8bit m2_597 (image2[91],filter_2[3],mul2_out[199][6]);
mul_20x8bit m2_598 (image2[92],filter_2[4],mul2_out[199][7]);
mul_20x8bit m2_599 (image2[93],filter_2[5],mul2_out[199][8]);
mul_20x8bit m2_600 (image2[104],filter_2[6],mul2_out[200][6]);
mul_20x8bit m2_601 (image2[105],filter_2[7],mul2_out[200][7]);
mul_20x8bit m2_602 (image2[106],filter_2[8],mul2_out[200][8]);

adder_24bit ad2_66 (mul2_out[198][6],mul2_out[198][7],mul2_out[198][8],mul2_out[199][6],mul2_out[199][7],mul2_out[199][8],mul2_out[200][6],mul2_out[200][7],mul2_out[200][8],conv2_out[66]);



mul_20x8bit m2_603 (image2[79],filter_2[0],mul2_out[201][6]);
mul_20x8bit m2_604 (image2[80],filter_2[1],mul2_out[201][7]);
mul_20x8bit m2_605 (image2[81],filter_2[2],mul2_out[201][8]);
mul_20x8bit m2_606 (image2[92],filter_2[3],mul2_out[202][6]);
mul_20x8bit m2_607 (image2[93],filter_2[4],mul2_out[202][7]);
mul_20x8bit m2_608 (image2[94],filter_2[5],mul2_out[202][8]);
mul_20x8bit m2_609 (image2[105],filter_2[6],mul2_out[203][6]);
mul_20x8bit m2_610 (image2[106],filter_2[7],mul2_out[203][7]);
mul_20x8bit m2_611 (image2[107],filter_2[8],mul2_out[203][8]);

adder_24bit ad2_67 (mul2_out[201][6],mul2_out[201][7],mul2_out[201][8],mul2_out[202][6],mul2_out[202][7],mul2_out[202][8],mul2_out[203][6],mul2_out[203][7],mul2_out[203][8],conv2_out[67]);



mul_20x8bit m2_612 (image2[80],filter_2[0],mul2_out[204][6]);
mul_20x8bit m2_613 (image2[81],filter_2[1],mul2_out[204][7]);
mul_20x8bit m2_614 (image2[82],filter_2[2],mul2_out[204][8]);
mul_20x8bit m2_615 (image2[93],filter_2[3],mul2_out[205][6]);
mul_20x8bit m2_616 (image2[94],filter_2[4],mul2_out[205][7]);
mul_20x8bit m2_617 (image2[95],filter_2[5],mul2_out[205][8]);
mul_20x8bit m2_618 (image2[106],filter_2[6],mul2_out[206][6]);
mul_20x8bit m2_619 (image2[107],filter_2[7],mul2_out[206][7]);
mul_20x8bit m2_620 (image2[108],filter_2[8],mul2_out[206][8]);

adder_24bit ad2_68 (mul2_out[204][6],mul2_out[204][7],mul2_out[204][8],mul2_out[205][6],mul2_out[205][7],mul2_out[205][8],mul2_out[206][6],mul2_out[206][7],mul2_out[206][8],conv2_out[68]);



mul_20x8bit m2_621 (image2[81],filter_2[0],mul2_out[207][6]);
mul_20x8bit m2_622 (image2[82],filter_2[1],mul2_out[207][7]);
mul_20x8bit m2_623 (image2[83],filter_2[2],mul2_out[207][8]);
mul_20x8bit m2_624 (image2[94],filter_2[3],mul2_out[208][6]);
mul_20x8bit m2_625 (image2[95],filter_2[4],mul2_out[208][7]);
mul_20x8bit m2_626 (image2[96],filter_2[5],mul2_out[208][8]);
mul_20x8bit m2_627 (image2[107],filter_2[6],mul2_out[209][6]);
mul_20x8bit m2_628 (image2[108],filter_2[7],mul2_out[209][7]);
mul_20x8bit m2_629 (image2[109],filter_2[8],mul2_out[209][8]);

adder_24bit ad2_69 (mul2_out[207][6],mul2_out[207][7],mul2_out[207][8],mul2_out[208][6],mul2_out[208][7],mul2_out[208][8],mul2_out[209][6],mul2_out[209][7],mul2_out[209][8],conv2_out[69]);



mul_20x8bit m2_630 (image2[82],filter_2[0],mul2_out[210][6]);
mul_20x8bit m2_631 (image2[83],filter_2[1],mul2_out[210][7]);
mul_20x8bit m2_632 (image2[84],filter_2[2],mul2_out[210][8]);
mul_20x8bit m2_633 (image2[95],filter_2[3],mul2_out[211][6]);
mul_20x8bit m2_634 (image2[96],filter_2[4],mul2_out[211][7]);
mul_20x8bit m2_635 (image2[97],filter_2[5],mul2_out[211][8]);
mul_20x8bit m2_636 (image2[108],filter_2[6],mul2_out[212][6]);
mul_20x8bit m2_637 (image2[109],filter_2[7],mul2_out[212][7]);
mul_20x8bit m2_638 (image2[110],filter_2[8],mul2_out[212][8]);

adder_24bit ad2_70 (mul2_out[210][6],mul2_out[210][7],mul2_out[210][8],mul2_out[211][6],mul2_out[211][7],mul2_out[211][8],mul2_out[212][6],mul2_out[212][7],mul2_out[212][8],conv2_out[70]);



mul_20x8bit m2_639 (image2[83],filter_2[0],mul2_out[213][6]);
mul_20x8bit m2_640 (image2[84],filter_2[1],mul2_out[213][7]);
mul_20x8bit m2_641 (image2[85],filter_2[2],mul2_out[213][8]);
mul_20x8bit m2_642 (image2[96],filter_2[3],mul2_out[214][6]);
mul_20x8bit m2_643 (image2[97],filter_2[4],mul2_out[214][7]);
mul_20x8bit m2_644 (image2[98],filter_2[5],mul2_out[214][8]);
mul_20x8bit m2_645 (image2[109],filter_2[6],mul2_out[215][6]);
mul_20x8bit m2_646 (image2[110],filter_2[7],mul2_out[215][7]);
mul_20x8bit m2_647 (image2[111],filter_2[8],mul2_out[215][8]);

adder_24bit ad2_71 (mul2_out[213][6],mul2_out[213][7],mul2_out[213][8],mul2_out[214][6],mul2_out[214][7],mul2_out[214][8],mul2_out[215][6],mul2_out[215][7],mul2_out[215][8],conv2_out[71]);



mul_20x8bit m2_648 (image2[84],filter_2[0],mul2_out[216][6]);
mul_20x8bit m2_649 (image2[85],filter_2[1],mul2_out[216][7]);
mul_20x8bit m2_650 (image2[86],filter_2[2],mul2_out[216][8]);
mul_20x8bit m2_651 (image2[97],filter_2[3],mul2_out[217][6]);
mul_20x8bit m2_652 (image2[98],filter_2[4],mul2_out[217][7]);
mul_20x8bit m2_653 (image2[99],filter_2[5],mul2_out[217][8]);
mul_20x8bit m2_654 (image2[110],filter_2[6],mul2_out[218][6]);
mul_20x8bit m2_655 (image2[111],filter_2[7],mul2_out[218][7]);
mul_20x8bit m2_656 (image2[112],filter_2[8],mul2_out[218][8]);

adder_24bit ad2_72 (mul2_out[216][6],mul2_out[216][7],mul2_out[216][8],mul2_out[217][6],mul2_out[217][7],mul2_out[217][8],mul2_out[218][6],mul2_out[218][7],mul2_out[218][8],conv2_out[72]);



mul_20x8bit m2_657 (image2[85],filter_2[0],mul2_out[219][6]);
mul_20x8bit m2_658 (image2[86],filter_2[1],mul2_out[219][7]);
mul_20x8bit m2_659 (image2[87],filter_2[2],mul2_out[219][8]);
mul_20x8bit m2_660 (image2[98],filter_2[3],mul2_out[220][6]);
mul_20x8bit m2_661 (image2[99],filter_2[4],mul2_out[220][7]);
mul_20x8bit m2_662 (image2[100],filter_2[5],mul2_out[220][8]);
mul_20x8bit m2_663 (image2[111],filter_2[6],mul2_out[221][6]);
mul_20x8bit m2_664 (image2[112],filter_2[7],mul2_out[221][7]);
mul_20x8bit m2_665 (image2[113],filter_2[8],mul2_out[221][8]);

adder_24bit ad2_73 (mul2_out[219][6],mul2_out[219][7],mul2_out[219][8],mul2_out[220][6],mul2_out[220][7],mul2_out[220][8],mul2_out[221][6],mul2_out[221][7],mul2_out[221][8],conv2_out[73]);



mul_20x8bit m2_666 (image2[86],filter_2[0],mul2_out[222][6]);
mul_20x8bit m2_667 (image2[87],filter_2[1],mul2_out[222][7]);
mul_20x8bit m2_668 (image2[88],filter_2[2],mul2_out[222][8]);
mul_20x8bit m2_669 (image2[99],filter_2[3],mul2_out[223][6]);
mul_20x8bit m2_670 (image2[100],filter_2[4],mul2_out[223][7]);
mul_20x8bit m2_671 (image2[101],filter_2[5],mul2_out[223][8]);
mul_20x8bit m2_672 (image2[112],filter_2[6],mul2_out[224][6]);
mul_20x8bit m2_673 (image2[113],filter_2[7],mul2_out[224][7]);
mul_20x8bit m2_674 (image2[114],filter_2[8],mul2_out[224][8]);

adder_24bit ad2_74 (mul2_out[222][6],mul2_out[222][7],mul2_out[222][8],mul2_out[223][6],mul2_out[223][7],mul2_out[223][8],mul2_out[224][6],mul2_out[224][7],mul2_out[224][8],conv2_out[74]);



mul_20x8bit m2_675 (image2[87],filter_2[0],mul2_out[225][6]);
mul_20x8bit m2_676 (image2[88],filter_2[1],mul2_out[225][7]);
mul_20x8bit m2_677 (image2[89],filter_2[2],mul2_out[225][8]);
mul_20x8bit m2_678 (image2[100],filter_2[3],mul2_out[226][6]);
mul_20x8bit m2_679 (image2[101],filter_2[4],mul2_out[226][7]);
mul_20x8bit m2_680 (image2[102],filter_2[5],mul2_out[226][8]);
mul_20x8bit m2_681 (image2[113],filter_2[6],mul2_out[227][6]);
mul_20x8bit m2_682 (image2[114],filter_2[7],mul2_out[227][7]);
mul_20x8bit m2_683 (image2[115],filter_2[8],mul2_out[227][8]);

adder_24bit ad2_75 (mul2_out[225][6],mul2_out[225][7],mul2_out[225][8],mul2_out[226][6],mul2_out[226][7],mul2_out[226][8],mul2_out[227][6],mul2_out[227][7],mul2_out[227][8],conv2_out[75]);



mul_20x8bit m2_684 (image2[88],filter_2[0],mul2_out[228][6]);
mul_20x8bit m2_685 (image2[89],filter_2[1],mul2_out[228][7]);
mul_20x8bit m2_686 (image2[90],filter_2[2],mul2_out[228][8]);
mul_20x8bit m2_687 (image2[101],filter_2[3],mul2_out[229][6]);
mul_20x8bit m2_688 (image2[102],filter_2[4],mul2_out[229][7]);
mul_20x8bit m2_689 (image2[103],filter_2[5],mul2_out[229][8]);
mul_20x8bit m2_690 (image2[114],filter_2[6],mul2_out[230][6]);
mul_20x8bit m2_691 (image2[115],filter_2[7],mul2_out[230][7]);
mul_20x8bit m2_692 (image2[116],filter_2[8],mul2_out[230][8]);

adder_24bit ad2_76 (mul2_out[228][6],mul2_out[228][7],mul2_out[228][8],mul2_out[229][6],mul2_out[229][7],mul2_out[229][8],mul2_out[230][6],mul2_out[230][7],mul2_out[230][8],conv2_out[76]);



mul_20x8bit m2_693 (image2[91],filter_2[0],mul2_out[231][7]);
mul_20x8bit m2_694 (image2[92],filter_2[1],mul2_out[231][8]);
mul_20x8bit m2_695 (image2[93],filter_2[2],mul2_out[231][9]);
mul_20x8bit m2_696 (image2[104],filter_2[3],mul2_out[232][7]);
mul_20x8bit m2_697 (image2[105],filter_2[4],mul2_out[232][8]);
mul_20x8bit m2_698 (image2[106],filter_2[5],mul2_out[232][9]);
mul_20x8bit m2_699 (image2[117],filter_2[6],mul2_out[233][7]);
mul_20x8bit m2_700 (image2[118],filter_2[7],mul2_out[233][8]);
mul_20x8bit m2_701 (image2[119],filter_2[8],mul2_out[233][9]);

adder_24bit ad2_77 (mul2_out[231][7],mul2_out[231][8],mul2_out[231][9],mul2_out[232][7],mul2_out[232][8],mul2_out[232][9],mul2_out[233][7],mul2_out[233][8],mul2_out[233][9],conv2_out[77]);



mul_20x8bit m2_702 (image2[92],filter_2[0],mul2_out[234][7]);
mul_20x8bit m2_703 (image2[93],filter_2[1],mul2_out[234][8]);
mul_20x8bit m2_704 (image2[94],filter_2[2],mul2_out[234][9]);
mul_20x8bit m2_705 (image2[105],filter_2[3],mul2_out[235][7]);
mul_20x8bit m2_706 (image2[106],filter_2[4],mul2_out[235][8]);
mul_20x8bit m2_707 (image2[107],filter_2[5],mul2_out[235][9]);
mul_20x8bit m2_708 (image2[118],filter_2[6],mul2_out[236][7]);
mul_20x8bit m2_709 (image2[119],filter_2[7],mul2_out[236][8]);
mul_20x8bit m2_710 (image2[120],filter_2[8],mul2_out[236][9]);

adder_24bit ad2_78 (mul2_out[234][7],mul2_out[234][8],mul2_out[234][9],mul2_out[235][7],mul2_out[235][8],mul2_out[235][9],mul2_out[236][7],mul2_out[236][8],mul2_out[236][9],conv2_out[78]);



mul_20x8bit m2_711 (image2[93],filter_2[0],mul2_out[237][7]);
mul_20x8bit m2_712 (image2[94],filter_2[1],mul2_out[237][8]);
mul_20x8bit m2_713 (image2[95],filter_2[2],mul2_out[237][9]);
mul_20x8bit m2_714 (image2[106],filter_2[3],mul2_out[238][7]);
mul_20x8bit m2_715 (image2[107],filter_2[4],mul2_out[238][8]);
mul_20x8bit m2_716 (image2[108],filter_2[5],mul2_out[238][9]);
mul_20x8bit m2_717 (image2[119],filter_2[6],mul2_out[239][7]);
mul_20x8bit m2_718 (image2[120],filter_2[7],mul2_out[239][8]);
mul_20x8bit m2_719 (image2[121],filter_2[8],mul2_out[239][9]);

adder_24bit ad2_79 (mul2_out[237][7],mul2_out[237][8],mul2_out[237][9],mul2_out[238][7],mul2_out[238][8],mul2_out[238][9],mul2_out[239][7],mul2_out[239][8],mul2_out[239][9],conv2_out[79]);



mul_20x8bit m2_720 (image2[94],filter_2[0],mul2_out[240][7]);
mul_20x8bit m2_721 (image2[95],filter_2[1],mul2_out[240][8]);
mul_20x8bit m2_722 (image2[96],filter_2[2],mul2_out[240][9]);
mul_20x8bit m2_723 (image2[107],filter_2[3],mul2_out[241][7]);
mul_20x8bit m2_724 (image2[108],filter_2[4],mul2_out[241][8]);
mul_20x8bit m2_725 (image2[109],filter_2[5],mul2_out[241][9]);
mul_20x8bit m2_726 (image2[120],filter_2[6],mul2_out[242][7]);
mul_20x8bit m2_727 (image2[121],filter_2[7],mul2_out[242][8]);
mul_20x8bit m2_728 (image2[122],filter_2[8],mul2_out[242][9]);

adder_24bit ad2_80 (mul2_out[240][7],mul2_out[240][8],mul2_out[240][9],mul2_out[241][7],mul2_out[241][8],mul2_out[241][9],mul2_out[242][7],mul2_out[242][8],mul2_out[242][9],conv2_out[80]);



mul_20x8bit m2_729 (image2[95],filter_2[0],mul2_out[243][7]);
mul_20x8bit m2_730 (image2[96],filter_2[1],mul2_out[243][8]);
mul_20x8bit m2_731 (image2[97],filter_2[2],mul2_out[243][9]);
mul_20x8bit m2_732 (image2[108],filter_2[3],mul2_out[244][7]);
mul_20x8bit m2_733 (image2[109],filter_2[4],mul2_out[244][8]);
mul_20x8bit m2_734 (image2[110],filter_2[5],mul2_out[244][9]);
mul_20x8bit m2_735 (image2[121],filter_2[6],mul2_out[245][7]);
mul_20x8bit m2_736 (image2[122],filter_2[7],mul2_out[245][8]);
mul_20x8bit m2_737 (image2[123],filter_2[8],mul2_out[245][9]);

adder_24bit ad2_81 (mul2_out[243][7],mul2_out[243][8],mul2_out[243][9],mul2_out[244][7],mul2_out[244][8],mul2_out[244][9],mul2_out[245][7],mul2_out[245][8],mul2_out[245][9],conv2_out[81]);



mul_20x8bit m2_738 (image2[96],filter_2[0],mul2_out[246][7]);
mul_20x8bit m2_739 (image2[97],filter_2[1],mul2_out[246][8]);
mul_20x8bit m2_740 (image2[98],filter_2[2],mul2_out[246][9]);
mul_20x8bit m2_741 (image2[109],filter_2[3],mul2_out[247][7]);
mul_20x8bit m2_742 (image2[110],filter_2[4],mul2_out[247][8]);
mul_20x8bit m2_743 (image2[111],filter_2[5],mul2_out[247][9]);
mul_20x8bit m2_744 (image2[122],filter_2[6],mul2_out[248][7]);
mul_20x8bit m2_745 (image2[123],filter_2[7],mul2_out[248][8]);
mul_20x8bit m2_746 (image2[124],filter_2[8],mul2_out[248][9]);

adder_24bit ad2_82 (mul2_out[246][7],mul2_out[246][8],mul2_out[246][9],mul2_out[247][7],mul2_out[247][8],mul2_out[247][9],mul2_out[248][7],mul2_out[248][8],mul2_out[248][9],conv2_out[82]);



mul_20x8bit m2_747 (image2[97],filter_2[0],mul2_out[249][7]);
mul_20x8bit m2_748 (image2[98],filter_2[1],mul2_out[249][8]);
mul_20x8bit m2_749 (image2[99],filter_2[2],mul2_out[249][9]);
mul_20x8bit m2_750 (image2[110],filter_2[3],mul2_out[250][7]);
mul_20x8bit m2_751 (image2[111],filter_2[4],mul2_out[250][8]);
mul_20x8bit m2_752 (image2[112],filter_2[5],mul2_out[250][9]);
mul_20x8bit m2_753 (image2[123],filter_2[6],mul2_out[251][7]);
mul_20x8bit m2_754 (image2[124],filter_2[7],mul2_out[251][8]);
mul_20x8bit m2_755 (image2[125],filter_2[8],mul2_out[251][9]);

adder_24bit ad2_83 (mul2_out[249][7],mul2_out[249][8],mul2_out[249][9],mul2_out[250][7],mul2_out[250][8],mul2_out[250][9],mul2_out[251][7],mul2_out[251][8],mul2_out[251][9],conv2_out[83]);



mul_20x8bit m2_756 (image2[98],filter_2[0],mul2_out[252][7]);
mul_20x8bit m2_757 (image2[99],filter_2[1],mul2_out[252][8]);
mul_20x8bit m2_758 (image2[100],filter_2[2],mul2_out[252][9]);
mul_20x8bit m2_759 (image2[111],filter_2[3],mul2_out[253][7]);
mul_20x8bit m2_760 (image2[112],filter_2[4],mul2_out[253][8]);
mul_20x8bit m2_761 (image2[113],filter_2[5],mul2_out[253][9]);
mul_20x8bit m2_762 (image2[124],filter_2[6],mul2_out[254][7]);
mul_20x8bit m2_763 (image2[125],filter_2[7],mul2_out[254][8]);
mul_20x8bit m2_764 (image2[126],filter_2[8],mul2_out[254][9]);

adder_24bit ad2_84 (mul2_out[252][7],mul2_out[252][8],mul2_out[252][9],mul2_out[253][7],mul2_out[253][8],mul2_out[253][9],mul2_out[254][7],mul2_out[254][8],mul2_out[254][9],conv2_out[84]);



mul_20x8bit m2_765 (image2[99],filter_2[0],mul2_out[255][7]);
mul_20x8bit m2_766 (image2[100],filter_2[1],mul2_out[255][8]);
mul_20x8bit m2_767 (image2[101],filter_2[2],mul2_out[255][9]);
mul_20x8bit m2_768 (image2[112],filter_2[3],mul2_out[256][7]);
mul_20x8bit m2_769 (image2[113],filter_2[4],mul2_out[256][8]);
mul_20x8bit m2_770 (image2[114],filter_2[5],mul2_out[256][9]);
mul_20x8bit m2_771 (image2[125],filter_2[6],mul2_out[257][7]);
mul_20x8bit m2_772 (image2[126],filter_2[7],mul2_out[257][8]);
mul_20x8bit m2_773 (image2[127],filter_2[8],mul2_out[257][9]);

adder_24bit ad2_85 (mul2_out[255][7],mul2_out[255][8],mul2_out[255][9],mul2_out[256][7],mul2_out[256][8],mul2_out[256][9],mul2_out[257][7],mul2_out[257][8],mul2_out[257][9],conv2_out[85]);



mul_20x8bit m2_774 (image2[100],filter_2[0],mul2_out[258][7]);
mul_20x8bit m2_775 (image2[101],filter_2[1],mul2_out[258][8]);
mul_20x8bit m2_776 (image2[102],filter_2[2],mul2_out[258][9]);
mul_20x8bit m2_777 (image2[113],filter_2[3],mul2_out[259][7]);
mul_20x8bit m2_778 (image2[114],filter_2[4],mul2_out[259][8]);
mul_20x8bit m2_779 (image2[115],filter_2[5],mul2_out[259][9]);
mul_20x8bit m2_780 (image2[126],filter_2[6],mul2_out[260][7]);
mul_20x8bit m2_781 (image2[127],filter_2[7],mul2_out[260][8]);
mul_20x8bit m2_782 (image2[128],filter_2[8],mul2_out[260][9]);

adder_24bit ad2_86 (mul2_out[258][7],mul2_out[258][8],mul2_out[258][9],mul2_out[259][7],mul2_out[259][8],mul2_out[259][9],mul2_out[260][7],mul2_out[260][8],mul2_out[260][9],conv2_out[86]);



mul_20x8bit m2_783 (image2[101],filter_2[0],mul2_out[261][7]);
mul_20x8bit m2_784 (image2[102],filter_2[1],mul2_out[261][8]);
mul_20x8bit m2_785 (image2[103],filter_2[2],mul2_out[261][9]);
mul_20x8bit m2_786 (image2[114],filter_2[3],mul2_out[262][7]);
mul_20x8bit m2_787 (image2[115],filter_2[4],mul2_out[262][8]);
mul_20x8bit m2_788 (image2[116],filter_2[5],mul2_out[262][9]);
mul_20x8bit m2_789 (image2[127],filter_2[6],mul2_out[263][7]);
mul_20x8bit m2_790 (image2[128],filter_2[7],mul2_out[263][8]);
mul_20x8bit m2_791 (image2[129],filter_2[8],mul2_out[263][9]);

adder_24bit ad2_87 (mul2_out[261][7],mul2_out[261][8],mul2_out[261][9],mul2_out[262][7],mul2_out[262][8],mul2_out[262][9],mul2_out[263][7],mul2_out[263][8],mul2_out[263][9],conv2_out[87]);



mul_20x8bit m2_792 (image2[104],filter_2[0],mul2_out[264][8]);
mul_20x8bit m2_793 (image2[105],filter_2[1],mul2_out[264][9]);
mul_20x8bit m2_794 (image2[106],filter_2[2],mul2_out[264][10]);
mul_20x8bit m2_795 (image2[117],filter_2[3],mul2_out[265][8]);
mul_20x8bit m2_796 (image2[118],filter_2[4],mul2_out[265][9]);
mul_20x8bit m2_797 (image2[119],filter_2[5],mul2_out[265][10]);
mul_20x8bit m2_798 (image2[130],filter_2[6],mul2_out[266][8]);
mul_20x8bit m2_799 (image2[131],filter_2[7],mul2_out[266][9]);
mul_20x8bit m2_800 (image2[132],filter_2[8],mul2_out[266][10]);

adder_24bit ad2_88 (mul2_out[264][8],mul2_out[264][9],mul2_out[264][10],mul2_out[265][8],mul2_out[265][9],mul2_out[265][10],mul2_out[266][8],mul2_out[266][9],mul2_out[266][10],conv2_out[88]);



mul_20x8bit m2_801 (image2[105],filter_2[0],mul2_out[267][8]);
mul_20x8bit m2_802 (image2[106],filter_2[1],mul2_out[267][9]);
mul_20x8bit m2_803 (image2[107],filter_2[2],mul2_out[267][10]);
mul_20x8bit m2_804 (image2[118],filter_2[3],mul2_out[268][8]);
mul_20x8bit m2_805 (image2[119],filter_2[4],mul2_out[268][9]);
mul_20x8bit m2_806 (image2[120],filter_2[5],mul2_out[268][10]);
mul_20x8bit m2_807 (image2[131],filter_2[6],mul2_out[269][8]);
mul_20x8bit m2_808 (image2[132],filter_2[7],mul2_out[269][9]);
mul_20x8bit m2_809 (image2[133],filter_2[8],mul2_out[269][10]);

adder_24bit ad2_89 (mul2_out[267][8],mul2_out[267][9],mul2_out[267][10],mul2_out[268][8],mul2_out[268][9],mul2_out[268][10],mul2_out[269][8],mul2_out[269][9],mul2_out[269][10],conv2_out[89]);



mul_20x8bit m2_810 (image2[106],filter_2[0],mul2_out[270][8]);
mul_20x8bit m2_811 (image2[107],filter_2[1],mul2_out[270][9]);
mul_20x8bit m2_812 (image2[108],filter_2[2],mul2_out[270][10]);
mul_20x8bit m2_813 (image2[119],filter_2[3],mul2_out[271][8]);
mul_20x8bit m2_814 (image2[120],filter_2[4],mul2_out[271][9]);
mul_20x8bit m2_815 (image2[121],filter_2[5],mul2_out[271][10]);
mul_20x8bit m2_816 (image2[132],filter_2[6],mul2_out[272][8]);
mul_20x8bit m2_817 (image2[133],filter_2[7],mul2_out[272][9]);
mul_20x8bit m2_818 (image2[134],filter_2[8],mul2_out[272][10]);

adder_24bit ad2_90 (mul2_out[270][8],mul2_out[270][9],mul2_out[270][10],mul2_out[271][8],mul2_out[271][9],mul2_out[271][10],mul2_out[272][8],mul2_out[272][9],mul2_out[272][10],conv2_out[90]);



mul_20x8bit m2_819 (image2[107],filter_2[0],mul2_out[273][8]);
mul_20x8bit m2_820 (image2[108],filter_2[1],mul2_out[273][9]);
mul_20x8bit m2_821 (image2[109],filter_2[2],mul2_out[273][10]);
mul_20x8bit m2_822 (image2[120],filter_2[3],mul2_out[274][8]);
mul_20x8bit m2_823 (image2[121],filter_2[4],mul2_out[274][9]);
mul_20x8bit m2_824 (image2[122],filter_2[5],mul2_out[274][10]);
mul_20x8bit m2_825 (image2[133],filter_2[6],mul2_out[275][8]);
mul_20x8bit m2_826 (image2[134],filter_2[7],mul2_out[275][9]);
mul_20x8bit m2_827 (image2[135],filter_2[8],mul2_out[275][10]);

adder_24bit ad2_91 (mul2_out[273][8],mul2_out[273][9],mul2_out[273][10],mul2_out[274][8],mul2_out[274][9],mul2_out[274][10],mul2_out[275][8],mul2_out[275][9],mul2_out[275][10],conv2_out[91]);



mul_20x8bit m2_828 (image2[108],filter_2[0],mul2_out[276][8]);
mul_20x8bit m2_829 (image2[109],filter_2[1],mul2_out[276][9]);
mul_20x8bit m2_830 (image2[110],filter_2[2],mul2_out[276][10]);
mul_20x8bit m2_831 (image2[121],filter_2[3],mul2_out[277][8]);
mul_20x8bit m2_832 (image2[122],filter_2[4],mul2_out[277][9]);
mul_20x8bit m2_833 (image2[123],filter_2[5],mul2_out[277][10]);
mul_20x8bit m2_834 (image2[134],filter_2[6],mul2_out[278][8]);
mul_20x8bit m2_835 (image2[135],filter_2[7],mul2_out[278][9]);
mul_20x8bit m2_836 (image2[136],filter_2[8],mul2_out[278][10]);

adder_24bit ad2_92 (mul2_out[276][8],mul2_out[276][9],mul2_out[276][10],mul2_out[277][8],mul2_out[277][9],mul2_out[277][10],mul2_out[278][8],mul2_out[278][9],mul2_out[278][10],conv2_out[92]);



mul_20x8bit m2_837 (image2[109],filter_2[0],mul2_out[279][8]);
mul_20x8bit m2_838 (image2[110],filter_2[1],mul2_out[279][9]);
mul_20x8bit m2_839 (image2[111],filter_2[2],mul2_out[279][10]);
mul_20x8bit m2_840 (image2[122],filter_2[3],mul2_out[280][8]);
mul_20x8bit m2_841 (image2[123],filter_2[4],mul2_out[280][9]);
mul_20x8bit m2_842 (image2[124],filter_2[5],mul2_out[280][10]);
mul_20x8bit m2_843 (image2[135],filter_2[6],mul2_out[281][8]);
mul_20x8bit m2_844 (image2[136],filter_2[7],mul2_out[281][9]);
mul_20x8bit m2_845 (image2[137],filter_2[8],mul2_out[281][10]);

adder_24bit ad2_93 (mul2_out[279][8],mul2_out[279][9],mul2_out[279][10],mul2_out[280][8],mul2_out[280][9],mul2_out[280][10],mul2_out[281][8],mul2_out[281][9],mul2_out[281][10],conv2_out[93]);



mul_20x8bit m2_846 (image2[110],filter_2[0],mul2_out[282][8]);
mul_20x8bit m2_847 (image2[111],filter_2[1],mul2_out[282][9]);
mul_20x8bit m2_848 (image2[112],filter_2[2],mul2_out[282][10]);
mul_20x8bit m2_849 (image2[123],filter_2[3],mul2_out[283][8]);
mul_20x8bit m2_850 (image2[124],filter_2[4],mul2_out[283][9]);
mul_20x8bit m2_851 (image2[125],filter_2[5],mul2_out[283][10]);
mul_20x8bit m2_852 (image2[136],filter_2[6],mul2_out[284][8]);
mul_20x8bit m2_853 (image2[137],filter_2[7],mul2_out[284][9]);
mul_20x8bit m2_854 (image2[138],filter_2[8],mul2_out[284][10]);

adder_24bit ad2_94 (mul2_out[282][8],mul2_out[282][9],mul2_out[282][10],mul2_out[283][8],mul2_out[283][9],mul2_out[283][10],mul2_out[284][8],mul2_out[284][9],mul2_out[284][10],conv2_out[94]);



mul_20x8bit m2_855 (image2[111],filter_2[0],mul2_out[285][8]);
mul_20x8bit m2_856 (image2[112],filter_2[1],mul2_out[285][9]);
mul_20x8bit m2_857 (image2[113],filter_2[2],mul2_out[285][10]);
mul_20x8bit m2_858 (image2[124],filter_2[3],mul2_out[286][8]);
mul_20x8bit m2_859 (image2[125],filter_2[4],mul2_out[286][9]);
mul_20x8bit m2_860 (image2[126],filter_2[5],mul2_out[286][10]);
mul_20x8bit m2_861 (image2[137],filter_2[6],mul2_out[287][8]);
mul_20x8bit m2_862 (image2[138],filter_2[7],mul2_out[287][9]);
mul_20x8bit m2_863 (image2[139],filter_2[8],mul2_out[287][10]);

adder_24bit ad2_95 (mul2_out[285][8],mul2_out[285][9],mul2_out[285][10],mul2_out[286][8],mul2_out[286][9],mul2_out[286][10],mul2_out[287][8],mul2_out[287][9],mul2_out[287][10],conv2_out[95]);



mul_20x8bit m2_864 (image2[112],filter_2[0],mul2_out[288][8]);
mul_20x8bit m2_865 (image2[113],filter_2[1],mul2_out[288][9]);
mul_20x8bit m2_866 (image2[114],filter_2[2],mul2_out[288][10]);
mul_20x8bit m2_867 (image2[125],filter_2[3],mul2_out[289][8]);
mul_20x8bit m2_868 (image2[126],filter_2[4],mul2_out[289][9]);
mul_20x8bit m2_869 (image2[127],filter_2[5],mul2_out[289][10]);
mul_20x8bit m2_870 (image2[138],filter_2[6],mul2_out[290][8]);
mul_20x8bit m2_871 (image2[139],filter_2[7],mul2_out[290][9]);
mul_20x8bit m2_872 (image2[140],filter_2[8],mul2_out[290][10]);

adder_24bit ad2_96 (mul2_out[288][8],mul2_out[288][9],mul2_out[288][10],mul2_out[289][8],mul2_out[289][9],mul2_out[289][10],mul2_out[290][8],mul2_out[290][9],mul2_out[290][10],conv2_out[96]);



mul_20x8bit m2_873 (image2[113],filter_2[0],mul2_out[291][8]);
mul_20x8bit m2_874 (image2[114],filter_2[1],mul2_out[291][9]);
mul_20x8bit m2_875 (image2[115],filter_2[2],mul2_out[291][10]);
mul_20x8bit m2_876 (image2[126],filter_2[3],mul2_out[292][8]);
mul_20x8bit m2_877 (image2[127],filter_2[4],mul2_out[292][9]);
mul_20x8bit m2_878 (image2[128],filter_2[5],mul2_out[292][10]);
mul_20x8bit m2_879 (image2[139],filter_2[6],mul2_out[293][8]);
mul_20x8bit m2_880 (image2[140],filter_2[7],mul2_out[293][9]);
mul_20x8bit m2_881 (image2[141],filter_2[8],mul2_out[293][10]);

adder_24bit ad2_97 (mul2_out[291][8],mul2_out[291][9],mul2_out[291][10],mul2_out[292][8],mul2_out[292][9],mul2_out[292][10],mul2_out[293][8],mul2_out[293][9],mul2_out[293][10],conv2_out[97]);



mul_20x8bit m2_882 (image2[114],filter_2[0],mul2_out[294][8]);
mul_20x8bit m2_883 (image2[115],filter_2[1],mul2_out[294][9]);
mul_20x8bit m2_884 (image2[116],filter_2[2],mul2_out[294][10]);
mul_20x8bit m2_885 (image2[127],filter_2[3],mul2_out[295][8]);
mul_20x8bit m2_886 (image2[128],filter_2[4],mul2_out[295][9]);
mul_20x8bit m2_887 (image2[129],filter_2[5],mul2_out[295][10]);
mul_20x8bit m2_888 (image2[140],filter_2[6],mul2_out[296][8]);
mul_20x8bit m2_889 (image2[141],filter_2[7],mul2_out[296][9]);
mul_20x8bit m2_890 (image2[142],filter_2[8],mul2_out[296][10]);

adder_24bit ad2_98 (mul2_out[294][8],mul2_out[294][9],mul2_out[294][10],mul2_out[295][8],mul2_out[295][9],mul2_out[295][10],mul2_out[296][8],mul2_out[296][9],mul2_out[296][10],conv2_out[98]);



mul_20x8bit m2_891 (image2[117],filter_2[0],mul2_out[297][9]);
mul_20x8bit m2_892 (image2[118],filter_2[1],mul2_out[297][10]);
mul_20x8bit m2_893 (image2[119],filter_2[2],mul2_out[297][11]);
mul_20x8bit m2_894 (image2[130],filter_2[3],mul2_out[298][9]);
mul_20x8bit m2_895 (image2[131],filter_2[4],mul2_out[298][10]);
mul_20x8bit m2_896 (image2[132],filter_2[5],mul2_out[298][11]);
mul_20x8bit m2_897 (image2[143],filter_2[6],mul2_out[299][9]);
mul_20x8bit m2_898 (image2[144],filter_2[7],mul2_out[299][10]);
mul_20x8bit m2_899 (image2[145],filter_2[8],mul2_out[299][11]);

adder_24bit ad2_99 (mul2_out[297][9],mul2_out[297][10],mul2_out[297][11],mul2_out[298][9],mul2_out[298][10],mul2_out[298][11],mul2_out[299][9],mul2_out[299][10],mul2_out[299][11],conv2_out[99]);



mul_20x8bit m2_900 (image2[118],filter_2[0],mul2_out[300][9]);
mul_20x8bit m2_901 (image2[119],filter_2[1],mul2_out[300][10]);
mul_20x8bit m2_902 (image2[120],filter_2[2],mul2_out[300][11]);
mul_20x8bit m2_903 (image2[131],filter_2[3],mul2_out[301][9]);
mul_20x8bit m2_904 (image2[132],filter_2[4],mul2_out[301][10]);
mul_20x8bit m2_905 (image2[133],filter_2[5],mul2_out[301][11]);
mul_20x8bit m2_906 (image2[144],filter_2[6],mul2_out[302][9]);
mul_20x8bit m2_907 (image2[145],filter_2[7],mul2_out[302][10]);
mul_20x8bit m2_908 (image2[146],filter_2[8],mul2_out[302][11]);

adder_24bit ad2_100 (mul2_out[300][9],mul2_out[300][10],mul2_out[300][11],mul2_out[301][9],mul2_out[301][10],mul2_out[301][11],mul2_out[302][9],mul2_out[302][10],mul2_out[302][11],conv2_out[100]);



mul_20x8bit m2_909 (image2[119],filter_2[0],mul2_out[303][9]);
mul_20x8bit m2_910 (image2[120],filter_2[1],mul2_out[303][10]);
mul_20x8bit m2_911 (image2[121],filter_2[2],mul2_out[303][11]);
mul_20x8bit m2_912 (image2[132],filter_2[3],mul2_out[304][9]);
mul_20x8bit m2_913 (image2[133],filter_2[4],mul2_out[304][10]);
mul_20x8bit m2_914 (image2[134],filter_2[5],mul2_out[304][11]);
mul_20x8bit m2_915 (image2[145],filter_2[6],mul2_out[305][9]);
mul_20x8bit m2_916 (image2[146],filter_2[7],mul2_out[305][10]);
mul_20x8bit m2_917 (image2[147],filter_2[8],mul2_out[305][11]);

adder_24bit ad2_101 (mul2_out[303][9],mul2_out[303][10],mul2_out[303][11],mul2_out[304][9],mul2_out[304][10],mul2_out[304][11],mul2_out[305][9],mul2_out[305][10],mul2_out[305][11],conv2_out[101]);



mul_20x8bit m2_918 (image2[120],filter_2[0],mul2_out[306][9]);
mul_20x8bit m2_919 (image2[121],filter_2[1],mul2_out[306][10]);
mul_20x8bit m2_920 (image2[122],filter_2[2],mul2_out[306][11]);
mul_20x8bit m2_921 (image2[133],filter_2[3],mul2_out[307][9]);
mul_20x8bit m2_922 (image2[134],filter_2[4],mul2_out[307][10]);
mul_20x8bit m2_923 (image2[135],filter_2[5],mul2_out[307][11]);
mul_20x8bit m2_924 (image2[146],filter_2[6],mul2_out[308][9]);
mul_20x8bit m2_925 (image2[147],filter_2[7],mul2_out[308][10]);
mul_20x8bit m2_926 (image2[148],filter_2[8],mul2_out[308][11]);

adder_24bit ad2_102 (mul2_out[306][9],mul2_out[306][10],mul2_out[306][11],mul2_out[307][9],mul2_out[307][10],mul2_out[307][11],mul2_out[308][9],mul2_out[308][10],mul2_out[308][11],conv2_out[102]);



mul_20x8bit m2_927 (image2[121],filter_2[0],mul2_out[309][9]);
mul_20x8bit m2_928 (image2[122],filter_2[1],mul2_out[309][10]);
mul_20x8bit m2_929 (image2[123],filter_2[2],mul2_out[309][11]);
mul_20x8bit m2_930 (image2[134],filter_2[3],mul2_out[310][9]);
mul_20x8bit m2_931 (image2[135],filter_2[4],mul2_out[310][10]);
mul_20x8bit m2_932 (image2[136],filter_2[5],mul2_out[310][11]);
mul_20x8bit m2_933 (image2[147],filter_2[6],mul2_out[311][9]);
mul_20x8bit m2_934 (image2[148],filter_2[7],mul2_out[311][10]);
mul_20x8bit m2_935 (image2[149],filter_2[8],mul2_out[311][11]);

adder_24bit ad2_103 (mul2_out[309][9],mul2_out[309][10],mul2_out[309][11],mul2_out[310][9],mul2_out[310][10],mul2_out[310][11],mul2_out[311][9],mul2_out[311][10],mul2_out[311][11],conv2_out[103]);



mul_20x8bit m2_936 (image2[122],filter_2[0],mul2_out[312][9]);
mul_20x8bit m2_937 (image2[123],filter_2[1],mul2_out[312][10]);
mul_20x8bit m2_938 (image2[124],filter_2[2],mul2_out[312][11]);
mul_20x8bit m2_939 (image2[135],filter_2[3],mul2_out[313][9]);
mul_20x8bit m2_940 (image2[136],filter_2[4],mul2_out[313][10]);
mul_20x8bit m2_941 (image2[137],filter_2[5],mul2_out[313][11]);
mul_20x8bit m2_942 (image2[148],filter_2[6],mul2_out[314][9]);
mul_20x8bit m2_943 (image2[149],filter_2[7],mul2_out[314][10]);
mul_20x8bit m2_944 (image2[150],filter_2[8],mul2_out[314][11]);

adder_24bit ad2_104 (mul2_out[312][9],mul2_out[312][10],mul2_out[312][11],mul2_out[313][9],mul2_out[313][10],mul2_out[313][11],mul2_out[314][9],mul2_out[314][10],mul2_out[314][11],conv2_out[104]);



mul_20x8bit m2_945 (image2[123],filter_2[0],mul2_out[315][9]);
mul_20x8bit m2_946 (image2[124],filter_2[1],mul2_out[315][10]);
mul_20x8bit m2_947 (image2[125],filter_2[2],mul2_out[315][11]);
mul_20x8bit m2_948 (image2[136],filter_2[3],mul2_out[316][9]);
mul_20x8bit m2_949 (image2[137],filter_2[4],mul2_out[316][10]);
mul_20x8bit m2_950 (image2[138],filter_2[5],mul2_out[316][11]);
mul_20x8bit m2_951 (image2[149],filter_2[6],mul2_out[317][9]);
mul_20x8bit m2_952 (image2[150],filter_2[7],mul2_out[317][10]);
mul_20x8bit m2_953 (image2[151],filter_2[8],mul2_out[317][11]);

adder_24bit ad2_105 (mul2_out[315][9],mul2_out[315][10],mul2_out[315][11],mul2_out[316][9],mul2_out[316][10],mul2_out[316][11],mul2_out[317][9],mul2_out[317][10],mul2_out[317][11],conv2_out[105]);



mul_20x8bit m2_954 (image2[124],filter_2[0],mul2_out[318][9]);
mul_20x8bit m2_955 (image2[125],filter_2[1],mul2_out[318][10]);
mul_20x8bit m2_956 (image2[126],filter_2[2],mul2_out[318][11]);
mul_20x8bit m2_957 (image2[137],filter_2[3],mul2_out[319][9]);
mul_20x8bit m2_958 (image2[138],filter_2[4],mul2_out[319][10]);
mul_20x8bit m2_959 (image2[139],filter_2[5],mul2_out[319][11]);
mul_20x8bit m2_960 (image2[150],filter_2[6],mul2_out[320][9]);
mul_20x8bit m2_961 (image2[151],filter_2[7],mul2_out[320][10]);
mul_20x8bit m2_962 (image2[152],filter_2[8],mul2_out[320][11]);

adder_24bit ad2_106 (mul2_out[318][9],mul2_out[318][10],mul2_out[318][11],mul2_out[319][9],mul2_out[319][10],mul2_out[319][11],mul2_out[320][9],mul2_out[320][10],mul2_out[320][11],conv2_out[106]);



mul_20x8bit m2_963 (image2[125],filter_2[0],mul2_out[321][9]);
mul_20x8bit m2_964 (image2[126],filter_2[1],mul2_out[321][10]);
mul_20x8bit m2_965 (image2[127],filter_2[2],mul2_out[321][11]);
mul_20x8bit m2_966 (image2[138],filter_2[3],mul2_out[322][9]);
mul_20x8bit m2_967 (image2[139],filter_2[4],mul2_out[322][10]);
mul_20x8bit m2_968 (image2[140],filter_2[5],mul2_out[322][11]);
mul_20x8bit m2_969 (image2[151],filter_2[6],mul2_out[323][9]);
mul_20x8bit m2_970 (image2[152],filter_2[7],mul2_out[323][10]);
mul_20x8bit m2_971 (image2[153],filter_2[8],mul2_out[323][11]);

adder_24bit ad2_107 (mul2_out[321][9],mul2_out[321][10],mul2_out[321][11],mul2_out[322][9],mul2_out[322][10],mul2_out[322][11],mul2_out[323][9],mul2_out[323][10],mul2_out[323][11],conv2_out[107]);



mul_20x8bit m2_972 (image2[126],filter_2[0],mul2_out[324][9]);
mul_20x8bit m2_973 (image2[127],filter_2[1],mul2_out[324][10]);
mul_20x8bit m2_974 (image2[128],filter_2[2],mul2_out[324][11]);
mul_20x8bit m2_975 (image2[139],filter_2[3],mul2_out[325][9]);
mul_20x8bit m2_976 (image2[140],filter_2[4],mul2_out[325][10]);
mul_20x8bit m2_977 (image2[141],filter_2[5],mul2_out[325][11]);
mul_20x8bit m2_978 (image2[152],filter_2[6],mul2_out[326][9]);
mul_20x8bit m2_979 (image2[153],filter_2[7],mul2_out[326][10]);
mul_20x8bit m2_980 (image2[154],filter_2[8],mul2_out[326][11]);

adder_24bit ad2_108 (mul2_out[324][9],mul2_out[324][10],mul2_out[324][11],mul2_out[325][9],mul2_out[325][10],mul2_out[325][11],mul2_out[326][9],mul2_out[326][10],mul2_out[326][11],conv2_out[108]);



mul_20x8bit m2_981 (image2[127],filter_2[0],mul2_out[327][9]);
mul_20x8bit m2_982 (image2[128],filter_2[1],mul2_out[327][10]);
mul_20x8bit m2_983 (image2[129],filter_2[2],mul2_out[327][11]);
mul_20x8bit m2_984 (image2[140],filter_2[3],mul2_out[328][9]);
mul_20x8bit m2_985 (image2[141],filter_2[4],mul2_out[328][10]);
mul_20x8bit m2_986 (image2[142],filter_2[5],mul2_out[328][11]);
mul_20x8bit m2_987 (image2[153],filter_2[6],mul2_out[329][9]);
mul_20x8bit m2_988 (image2[154],filter_2[7],mul2_out[329][10]);
mul_20x8bit m2_989 (image2[155],filter_2[8],mul2_out[329][11]);

adder_24bit ad2_109 (mul2_out[327][9],mul2_out[327][10],mul2_out[327][11],mul2_out[328][9],mul2_out[328][10],mul2_out[328][11],mul2_out[329][9],mul2_out[329][10],mul2_out[329][11],conv2_out[109]);



mul_20x8bit m2_990 (image2[130],filter_2[0],mul2_out[330][10]);
mul_20x8bit m2_991 (image2[131],filter_2[1],mul2_out[330][11]);
mul_20x8bit m2_992 (image2[132],filter_2[2],mul2_out[330][12]);
mul_20x8bit m2_993 (image2[143],filter_2[3],mul2_out[331][10]);
mul_20x8bit m2_994 (image2[144],filter_2[4],mul2_out[331][11]);
mul_20x8bit m2_995 (image2[145],filter_2[5],mul2_out[331][12]);
mul_20x8bit m2_996 (image2[156],filter_2[6],mul2_out[332][10]);
mul_20x8bit m2_997 (image2[157],filter_2[7],mul2_out[332][11]);
mul_20x8bit m2_998 (image2[158],filter_2[8],mul2_out[332][12]);

adder_24bit ad2_110 (mul2_out[330][10],mul2_out[330][11],mul2_out[330][12],mul2_out[331][10],mul2_out[331][11],mul2_out[331][12],mul2_out[332][10],mul2_out[332][11],mul2_out[332][12],conv2_out[110]);



mul_20x8bit m2_999 (image2[131],filter_2[0],mul2_out[333][10]);
mul_20x8bit m2_1000 (image2[132],filter_2[1],mul2_out[333][11]);
mul_20x8bit m2_1001 (image2[133],filter_2[2],mul2_out[333][12]);
mul_20x8bit m2_1002 (image2[144],filter_2[3],mul2_out[334][10]);
mul_20x8bit m2_1003 (image2[145],filter_2[4],mul2_out[334][11]);
mul_20x8bit m2_1004 (image2[146],filter_2[5],mul2_out[334][12]);
mul_20x8bit m2_1005 (image2[157],filter_2[6],mul2_out[335][10]);
mul_20x8bit m2_1006 (image2[158],filter_2[7],mul2_out[335][11]);
mul_20x8bit m2_1007 (image2[159],filter_2[8],mul2_out[335][12]);

adder_24bit ad2_111 (mul2_out[333][10],mul2_out[333][11],mul2_out[333][12],mul2_out[334][10],mul2_out[334][11],mul2_out[334][12],mul2_out[335][10],mul2_out[335][11],mul2_out[335][12],conv2_out[111]);



mul_20x8bit m2_1008 (image2[132],filter_2[0],mul2_out[336][10]);
mul_20x8bit m2_1009 (image2[133],filter_2[1],mul2_out[336][11]);
mul_20x8bit m2_1010 (image2[134],filter_2[2],mul2_out[336][12]);
mul_20x8bit m2_1011 (image2[145],filter_2[3],mul2_out[337][10]);
mul_20x8bit m2_1012 (image2[146],filter_2[4],mul2_out[337][11]);
mul_20x8bit m2_1013 (image2[147],filter_2[5],mul2_out[337][12]);
mul_20x8bit m2_1014 (image2[158],filter_2[6],mul2_out[338][10]);
mul_20x8bit m2_1015 (image2[159],filter_2[7],mul2_out[338][11]);
mul_20x8bit m2_1016 (image2[160],filter_2[8],mul2_out[338][12]);

adder_24bit ad2_112 (mul2_out[336][10],mul2_out[336][11],mul2_out[336][12],mul2_out[337][10],mul2_out[337][11],mul2_out[337][12],mul2_out[338][10],mul2_out[338][11],mul2_out[338][12],conv2_out[112]);



mul_20x8bit m2_1017 (image2[133],filter_2[0],mul2_out[339][10]);
mul_20x8bit m2_1018 (image2[134],filter_2[1],mul2_out[339][11]);
mul_20x8bit m2_1019 (image2[135],filter_2[2],mul2_out[339][12]);
mul_20x8bit m2_1020 (image2[146],filter_2[3],mul2_out[340][10]);
mul_20x8bit m2_1021 (image2[147],filter_2[4],mul2_out[340][11]);
mul_20x8bit m2_1022 (image2[148],filter_2[5],mul2_out[340][12]);
mul_20x8bit m2_1023 (image2[159],filter_2[6],mul2_out[341][10]);
mul_20x8bit m2_1024 (image2[160],filter_2[7],mul2_out[341][11]);
mul_20x8bit m2_1025 (image2[161],filter_2[8],mul2_out[341][12]);

adder_24bit ad2_113 (mul2_out[339][10],mul2_out[339][11],mul2_out[339][12],mul2_out[340][10],mul2_out[340][11],mul2_out[340][12],mul2_out[341][10],mul2_out[341][11],mul2_out[341][12],conv2_out[113]);



mul_20x8bit m2_1026 (image2[134],filter_2[0],mul2_out[342][10]);
mul_20x8bit m2_1027 (image2[135],filter_2[1],mul2_out[342][11]);
mul_20x8bit m2_1028 (image2[136],filter_2[2],mul2_out[342][12]);
mul_20x8bit m2_1029 (image2[147],filter_2[3],mul2_out[343][10]);
mul_20x8bit m2_1030 (image2[148],filter_2[4],mul2_out[343][11]);
mul_20x8bit m2_1031 (image2[149],filter_2[5],mul2_out[343][12]);
mul_20x8bit m2_1032 (image2[160],filter_2[6],mul2_out[344][10]);
mul_20x8bit m2_1033 (image2[161],filter_2[7],mul2_out[344][11]);
mul_20x8bit m2_1034 (image2[162],filter_2[8],mul2_out[344][12]);

adder_24bit ad2_114 (mul2_out[342][10],mul2_out[342][11],mul2_out[342][12],mul2_out[343][10],mul2_out[343][11],mul2_out[343][12],mul2_out[344][10],mul2_out[344][11],mul2_out[344][12],conv2_out[114]);



mul_20x8bit m2_1035 (image2[135],filter_2[0],mul2_out[345][10]);
mul_20x8bit m2_1036 (image2[136],filter_2[1],mul2_out[345][11]);
mul_20x8bit m2_1037 (image2[137],filter_2[2],mul2_out[345][12]);
mul_20x8bit m2_1038 (image2[148],filter_2[3],mul2_out[346][10]);
mul_20x8bit m2_1039 (image2[149],filter_2[4],mul2_out[346][11]);
mul_20x8bit m2_1040 (image2[150],filter_2[5],mul2_out[346][12]);
mul_20x8bit m2_1041 (image2[161],filter_2[6],mul2_out[347][10]);
mul_20x8bit m2_1042 (image2[162],filter_2[7],mul2_out[347][11]);
mul_20x8bit m2_1043 (image2[163],filter_2[8],mul2_out[347][12]);

adder_24bit ad2_115 (mul2_out[345][10],mul2_out[345][11],mul2_out[345][12],mul2_out[346][10],mul2_out[346][11],mul2_out[346][12],mul2_out[347][10],mul2_out[347][11],mul2_out[347][12],conv2_out[115]);



mul_20x8bit m2_1044 (image2[136],filter_2[0],mul2_out[348][10]);
mul_20x8bit m2_1045 (image2[137],filter_2[1],mul2_out[348][11]);
mul_20x8bit m2_1046 (image2[138],filter_2[2],mul2_out[348][12]);
mul_20x8bit m2_1047 (image2[149],filter_2[3],mul2_out[349][10]);
mul_20x8bit m2_1048 (image2[150],filter_2[4],mul2_out[349][11]);
mul_20x8bit m2_1049 (image2[151],filter_2[5],mul2_out[349][12]);
mul_20x8bit m2_1050 (image2[162],filter_2[6],mul2_out[350][10]);
mul_20x8bit m2_1051 (image2[163],filter_2[7],mul2_out[350][11]);
mul_20x8bit m2_1052 (image2[164],filter_2[8],mul2_out[350][12]);

adder_24bit ad2_116 (mul2_out[348][10],mul2_out[348][11],mul2_out[348][12],mul2_out[349][10],mul2_out[349][11],mul2_out[349][12],mul2_out[350][10],mul2_out[350][11],mul2_out[350][12],conv2_out[116]);



mul_20x8bit m2_1053 (image2[137],filter_2[0],mul2_out[351][10]);
mul_20x8bit m2_1054 (image2[138],filter_2[1],mul2_out[351][11]);
mul_20x8bit m2_1055 (image2[139],filter_2[2],mul2_out[351][12]);
mul_20x8bit m2_1056 (image2[150],filter_2[3],mul2_out[352][10]);
mul_20x8bit m2_1057 (image2[151],filter_2[4],mul2_out[352][11]);
mul_20x8bit m2_1058 (image2[152],filter_2[5],mul2_out[352][12]);
mul_20x8bit m2_1059 (image2[163],filter_2[6],mul2_out[353][10]);
mul_20x8bit m2_1060 (image2[164],filter_2[7],mul2_out[353][11]);
mul_20x8bit m2_1061 (image2[165],filter_2[8],mul2_out[353][12]);

adder_24bit ad2_117 (mul2_out[351][10],mul2_out[351][11],mul2_out[351][12],mul2_out[352][10],mul2_out[352][11],mul2_out[352][12],mul2_out[353][10],mul2_out[353][11],mul2_out[353][12],conv2_out[117]);



mul_20x8bit m2_1062 (image2[138],filter_2[0],mul2_out[354][10]);
mul_20x8bit m2_1063 (image2[139],filter_2[1],mul2_out[354][11]);
mul_20x8bit m2_1064 (image2[140],filter_2[2],mul2_out[354][12]);
mul_20x8bit m2_1065 (image2[151],filter_2[3],mul2_out[355][10]);
mul_20x8bit m2_1066 (image2[152],filter_2[4],mul2_out[355][11]);
mul_20x8bit m2_1067 (image2[153],filter_2[5],mul2_out[355][12]);
mul_20x8bit m2_1068 (image2[164],filter_2[6],mul2_out[356][10]);
mul_20x8bit m2_1069 (image2[165],filter_2[7],mul2_out[356][11]);
mul_20x8bit m2_1070 (image2[166],filter_2[8],mul2_out[356][12]);

adder_24bit ad2_118 (mul2_out[354][10],mul2_out[354][11],mul2_out[354][12],mul2_out[355][10],mul2_out[355][11],mul2_out[355][12],mul2_out[356][10],mul2_out[356][11],mul2_out[356][12],conv2_out[118]);



mul_20x8bit m2_1071 (image2[139],filter_2[0],mul2_out[357][10]);
mul_20x8bit m2_1072 (image2[140],filter_2[1],mul2_out[357][11]);
mul_20x8bit m2_1073 (image2[141],filter_2[2],mul2_out[357][12]);
mul_20x8bit m2_1074 (image2[152],filter_2[3],mul2_out[358][10]);
mul_20x8bit m2_1075 (image2[153],filter_2[4],mul2_out[358][11]);
mul_20x8bit m2_1076 (image2[154],filter_2[5],mul2_out[358][12]);
mul_20x8bit m2_1077 (image2[165],filter_2[6],mul2_out[359][10]);
mul_20x8bit m2_1078 (image2[166],filter_2[7],mul2_out[359][11]);
mul_20x8bit m2_1079 (image2[167],filter_2[8],mul2_out[359][12]);

adder_24bit ad2_119 (mul2_out[357][10],mul2_out[357][11],mul2_out[357][12],mul2_out[358][10],mul2_out[358][11],mul2_out[358][12],mul2_out[359][10],mul2_out[359][11],mul2_out[359][12],conv2_out[119]);



mul_20x8bit m2_1080 (image2[140],filter_2[0],mul2_out[360][10]);
mul_20x8bit m2_1081 (image2[141],filter_2[1],mul2_out[360][11]);
mul_20x8bit m2_1082 (image2[142],filter_2[2],mul2_out[360][12]);
mul_20x8bit m2_1083 (image2[153],filter_2[3],mul2_out[361][10]);
mul_20x8bit m2_1084 (image2[154],filter_2[4],mul2_out[361][11]);
mul_20x8bit m2_1085 (image2[155],filter_2[5],mul2_out[361][12]);
mul_20x8bit m2_1086 (image2[166],filter_2[6],mul2_out[362][10]);
mul_20x8bit m2_1087 (image2[167],filter_2[7],mul2_out[362][11]);
mul_20x8bit m2_1088 (image2[168],filter_2[8],mul2_out[362][12]);

adder_24bit ad2_120 (mul2_out[360][10],mul2_out[360][11],mul2_out[360][12],mul2_out[361][10],mul2_out[361][11],mul2_out[361][12],mul2_out[362][10],mul2_out[362][11],mul2_out[362][12],conv2_out[120]);
endmodule
