`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/10/2025 10:42:35 AM
// Design Name: 
// Module Name: CNN_conv1_final_mod
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module adder_8bit ( // with sign
input logic signed [15:0]a,b,c,d,e,f,g,h,hi,
output logic signed [19:0] sum //signed
);

assign sum = a+b+c+d+e+f+g+h+hi; // add all without sign bit
endmodule


module mul_8x8bit(
input logic signed [8:0]al, // 8bit a without signed and 8 bit 256
input logic signed [7:0]bl, // max number after mul with 256 is 63(6bit)7 bit with sign
output logic signed [15:0] mult_out
);

assign mult_out = al*bl; // multiply all without sign bit al[7:0]*bl[5:0]
endmodule


 module CNN_conv1_final_mod(
input logic clk,rst,
input logic signed [8:0] image[0:783], // unsigned
input logic signed [7:0]filter[0:8], // signed(max:63) kernel_1_re[4]3][3]: kernel_1_re[0][x][y],kernel_1_re[1][x][y], . kernel_1_re[3][x][y], round off 3 decimal points
output logic signed [19:0] conv_out [0:675] // signed
);
 logic signed [15:0] mul_out [0:2027][0:27]; // signed


mul_8x8bit m0 (image[0],filter[0],mul_out[0][0]);
mul_8x8bit m1 (image[1],filter[1],mul_out[0][1]);
mul_8x8bit m2 (image[2],filter[2],mul_out[0][2]);
mul_8x8bit m3 (image[28],filter[3],mul_out[1][0]);
mul_8x8bit m4 (image[29],filter[4],mul_out[1][1]);
mul_8x8bit m5 (image[30],filter[5],mul_out[1][2]);
mul_8x8bit m6 (image[56],filter[6],mul_out[2][0]);
mul_8x8bit m7 (image[57],filter[7],mul_out[2][1]);
mul_8x8bit m8 (image[58],filter[8],mul_out[2][2]);

adder_8bit ad0 (mul_out[0][0],mul_out[0][1],mul_out[0][2],mul_out[1][0],mul_out[1][1],mul_out[1][2],mul_out[2][0],mul_out[2][1],mul_out[2][2],conv_out[0]);



mul_8x8bit m9 (image[1],filter[0],mul_out[3][0]);
mul_8x8bit m10 (image[2],filter[1],mul_out[3][1]);
mul_8x8bit m11 (image[3],filter[2],mul_out[3][2]);
mul_8x8bit m12 (image[29],filter[3],mul_out[4][0]);
mul_8x8bit m13 (image[30],filter[4],mul_out[4][1]);
mul_8x8bit m14 (image[31],filter[5],mul_out[4][2]);
mul_8x8bit m15 (image[57],filter[6],mul_out[5][0]);
mul_8x8bit m16 (image[58],filter[7],mul_out[5][1]);
mul_8x8bit m17 (image[59],filter[8],mul_out[5][2]);

adder_8bit ad1 (mul_out[3][0],mul_out[3][1],mul_out[3][2],mul_out[4][0],mul_out[4][1],mul_out[4][2],mul_out[5][0],mul_out[5][1],mul_out[5][2],conv_out[1]);



mul_8x8bit m18 (image[2],filter[0],mul_out[6][0]);
mul_8x8bit m19 (image[3],filter[1],mul_out[6][1]);
mul_8x8bit m20 (image[4],filter[2],mul_out[6][2]);
mul_8x8bit m21 (image[30],filter[3],mul_out[7][0]);
mul_8x8bit m22 (image[31],filter[4],mul_out[7][1]);
mul_8x8bit m23 (image[32],filter[5],mul_out[7][2]);
mul_8x8bit m24 (image[58],filter[6],mul_out[8][0]);
mul_8x8bit m25 (image[59],filter[7],mul_out[8][1]);
mul_8x8bit m26 (image[60],filter[8],mul_out[8][2]);

adder_8bit ad2 (mul_out[6][0],mul_out[6][1],mul_out[6][2],mul_out[7][0],mul_out[7][1],mul_out[7][2],mul_out[8][0],mul_out[8][1],mul_out[8][2],conv_out[2]);



mul_8x8bit m27 (image[3],filter[0],mul_out[9][0]);
mul_8x8bit m28 (image[4],filter[1],mul_out[9][1]);
mul_8x8bit m29 (image[5],filter[2],mul_out[9][2]);
mul_8x8bit m30 (image[31],filter[3],mul_out[10][0]);
mul_8x8bit m31 (image[32],filter[4],mul_out[10][1]);
mul_8x8bit m32 (image[33],filter[5],mul_out[10][2]);
mul_8x8bit m33 (image[59],filter[6],mul_out[11][0]);
mul_8x8bit m34 (image[60],filter[7],mul_out[11][1]);
mul_8x8bit m35 (image[61],filter[8],mul_out[11][2]);

adder_8bit ad3 (mul_out[9][0],mul_out[9][1],mul_out[9][2],mul_out[10][0],mul_out[10][1],mul_out[10][2],mul_out[11][0],mul_out[11][1],mul_out[11][2],conv_out[3]);



mul_8x8bit m36 (image[4],filter[0],mul_out[12][0]);
mul_8x8bit m37 (image[5],filter[1],mul_out[12][1]);
mul_8x8bit m38 (image[6],filter[2],mul_out[12][2]);
mul_8x8bit m39 (image[32],filter[3],mul_out[13][0]);
mul_8x8bit m40 (image[33],filter[4],mul_out[13][1]);
mul_8x8bit m41 (image[34],filter[5],mul_out[13][2]);
mul_8x8bit m42 (image[60],filter[6],mul_out[14][0]);
mul_8x8bit m43 (image[61],filter[7],mul_out[14][1]);
mul_8x8bit m44 (image[62],filter[8],mul_out[14][2]);

adder_8bit ad4 (mul_out[12][0],mul_out[12][1],mul_out[12][2],mul_out[13][0],mul_out[13][1],mul_out[13][2],mul_out[14][0],mul_out[14][1],mul_out[14][2],conv_out[4]);



mul_8x8bit m45 (image[5],filter[0],mul_out[15][0]);
mul_8x8bit m46 (image[6],filter[1],mul_out[15][1]);
mul_8x8bit m47 (image[7],filter[2],mul_out[15][2]);
mul_8x8bit m48 (image[33],filter[3],mul_out[16][0]);
mul_8x8bit m49 (image[34],filter[4],mul_out[16][1]);
mul_8x8bit m50 (image[35],filter[5],mul_out[16][2]);
mul_8x8bit m51 (image[61],filter[6],mul_out[17][0]);
mul_8x8bit m52 (image[62],filter[7],mul_out[17][1]);
mul_8x8bit m53 (image[63],filter[8],mul_out[17][2]);

adder_8bit ad5 (mul_out[15][0],mul_out[15][1],mul_out[15][2],mul_out[16][0],mul_out[16][1],mul_out[16][2],mul_out[17][0],mul_out[17][1],mul_out[17][2],conv_out[5]);



mul_8x8bit m54 (image[6],filter[0],mul_out[18][0]);
mul_8x8bit m55 (image[7],filter[1],mul_out[18][1]);
mul_8x8bit m56 (image[8],filter[2],mul_out[18][2]);
mul_8x8bit m57 (image[34],filter[3],mul_out[19][0]);
mul_8x8bit m58 (image[35],filter[4],mul_out[19][1]);
mul_8x8bit m59 (image[36],filter[5],mul_out[19][2]);
mul_8x8bit m60 (image[62],filter[6],mul_out[20][0]);
mul_8x8bit m61 (image[63],filter[7],mul_out[20][1]);
mul_8x8bit m62 (image[64],filter[8],mul_out[20][2]);

adder_8bit ad6 (mul_out[18][0],mul_out[18][1],mul_out[18][2],mul_out[19][0],mul_out[19][1],mul_out[19][2],mul_out[20][0],mul_out[20][1],mul_out[20][2],conv_out[6]);



mul_8x8bit m63 (image[7],filter[0],mul_out[21][0]);
mul_8x8bit m64 (image[8],filter[1],mul_out[21][1]);
mul_8x8bit m65 (image[9],filter[2],mul_out[21][2]);
mul_8x8bit m66 (image[35],filter[3],mul_out[22][0]);
mul_8x8bit m67 (image[36],filter[4],mul_out[22][1]);
mul_8x8bit m68 (image[37],filter[5],mul_out[22][2]);
mul_8x8bit m69 (image[63],filter[6],mul_out[23][0]);
mul_8x8bit m70 (image[64],filter[7],mul_out[23][1]);
mul_8x8bit m71 (image[65],filter[8],mul_out[23][2]);

adder_8bit ad7 (mul_out[21][0],mul_out[21][1],mul_out[21][2],mul_out[22][0],mul_out[22][1],mul_out[22][2],mul_out[23][0],mul_out[23][1],mul_out[23][2],conv_out[7]);



mul_8x8bit m72 (image[8],filter[0],mul_out[24][0]);
mul_8x8bit m73 (image[9],filter[1],mul_out[24][1]);
mul_8x8bit m74 (image[10],filter[2],mul_out[24][2]);
mul_8x8bit m75 (image[36],filter[3],mul_out[25][0]);
mul_8x8bit m76 (image[37],filter[4],mul_out[25][1]);
mul_8x8bit m77 (image[38],filter[5],mul_out[25][2]);
mul_8x8bit m78 (image[64],filter[6],mul_out[26][0]);
mul_8x8bit m79 (image[65],filter[7],mul_out[26][1]);
mul_8x8bit m80 (image[66],filter[8],mul_out[26][2]);

adder_8bit ad8 (mul_out[24][0],mul_out[24][1],mul_out[24][2],mul_out[25][0],mul_out[25][1],mul_out[25][2],mul_out[26][0],mul_out[26][1],mul_out[26][2],conv_out[8]);



mul_8x8bit m81 (image[9],filter[0],mul_out[27][0]);
mul_8x8bit m82 (image[10],filter[1],mul_out[27][1]);
mul_8x8bit m83 (image[11],filter[2],mul_out[27][2]);
mul_8x8bit m84 (image[37],filter[3],mul_out[28][0]);
mul_8x8bit m85 (image[38],filter[4],mul_out[28][1]);
mul_8x8bit m86 (image[39],filter[5],mul_out[28][2]);
mul_8x8bit m87 (image[65],filter[6],mul_out[29][0]);
mul_8x8bit m88 (image[66],filter[7],mul_out[29][1]);
mul_8x8bit m89 (image[67],filter[8],mul_out[29][2]);

adder_8bit ad9 (mul_out[27][0],mul_out[27][1],mul_out[27][2],mul_out[28][0],mul_out[28][1],mul_out[28][2],mul_out[29][0],mul_out[29][1],mul_out[29][2],conv_out[9]);



mul_8x8bit m90 (image[10],filter[0],mul_out[30][0]);
mul_8x8bit m91 (image[11],filter[1],mul_out[30][1]);
mul_8x8bit m92 (image[12],filter[2],mul_out[30][2]);
mul_8x8bit m93 (image[38],filter[3],mul_out[31][0]);
mul_8x8bit m94 (image[39],filter[4],mul_out[31][1]);
mul_8x8bit m95 (image[40],filter[5],mul_out[31][2]);
mul_8x8bit m96 (image[66],filter[6],mul_out[32][0]);
mul_8x8bit m97 (image[67],filter[7],mul_out[32][1]);
mul_8x8bit m98 (image[68],filter[8],mul_out[32][2]);

adder_8bit ad10 (mul_out[30][0],mul_out[30][1],mul_out[30][2],mul_out[31][0],mul_out[31][1],mul_out[31][2],mul_out[32][0],mul_out[32][1],mul_out[32][2],conv_out[10]);



mul_8x8bit m99 (image[11],filter[0],mul_out[33][0]);
mul_8x8bit m100 (image[12],filter[1],mul_out[33][1]);
mul_8x8bit m101 (image[13],filter[2],mul_out[33][2]);
mul_8x8bit m102 (image[39],filter[3],mul_out[34][0]);
mul_8x8bit m103 (image[40],filter[4],mul_out[34][1]);
mul_8x8bit m104 (image[41],filter[5],mul_out[34][2]);
mul_8x8bit m105 (image[67],filter[6],mul_out[35][0]);
mul_8x8bit m106 (image[68],filter[7],mul_out[35][1]);
mul_8x8bit m107 (image[69],filter[8],mul_out[35][2]);

adder_8bit ad11 (mul_out[33][0],mul_out[33][1],mul_out[33][2],mul_out[34][0],mul_out[34][1],mul_out[34][2],mul_out[35][0],mul_out[35][1],mul_out[35][2],conv_out[11]);



mul_8x8bit m108 (image[12],filter[0],mul_out[36][0]);
mul_8x8bit m109 (image[13],filter[1],mul_out[36][1]);
mul_8x8bit m110 (image[14],filter[2],mul_out[36][2]);
mul_8x8bit m111 (image[40],filter[3],mul_out[37][0]);
mul_8x8bit m112 (image[41],filter[4],mul_out[37][1]);
mul_8x8bit m113 (image[42],filter[5],mul_out[37][2]);
mul_8x8bit m114 (image[68],filter[6],mul_out[38][0]);
mul_8x8bit m115 (image[69],filter[7],mul_out[38][1]);
mul_8x8bit m116 (image[70],filter[8],mul_out[38][2]);

adder_8bit ad12 (mul_out[36][0],mul_out[36][1],mul_out[36][2],mul_out[37][0],mul_out[37][1],mul_out[37][2],mul_out[38][0],mul_out[38][1],mul_out[38][2],conv_out[12]);



mul_8x8bit m117 (image[13],filter[0],mul_out[39][0]);
mul_8x8bit m118 (image[14],filter[1],mul_out[39][1]);
mul_8x8bit m119 (image[15],filter[2],mul_out[39][2]);
mul_8x8bit m120 (image[41],filter[3],mul_out[40][0]);
mul_8x8bit m121 (image[42],filter[4],mul_out[40][1]);
mul_8x8bit m122 (image[43],filter[5],mul_out[40][2]);
mul_8x8bit m123 (image[69],filter[6],mul_out[41][0]);
mul_8x8bit m124 (image[70],filter[7],mul_out[41][1]);
mul_8x8bit m125 (image[71],filter[8],mul_out[41][2]);

adder_8bit ad13 (mul_out[39][0],mul_out[39][1],mul_out[39][2],mul_out[40][0],mul_out[40][1],mul_out[40][2],mul_out[41][0],mul_out[41][1],mul_out[41][2],conv_out[13]);



mul_8x8bit m126 (image[14],filter[0],mul_out[42][0]);
mul_8x8bit m127 (image[15],filter[1],mul_out[42][1]);
mul_8x8bit m128 (image[16],filter[2],mul_out[42][2]);
mul_8x8bit m129 (image[42],filter[3],mul_out[43][0]);
mul_8x8bit m130 (image[43],filter[4],mul_out[43][1]);
mul_8x8bit m131 (image[44],filter[5],mul_out[43][2]);
mul_8x8bit m132 (image[70],filter[6],mul_out[44][0]);
mul_8x8bit m133 (image[71],filter[7],mul_out[44][1]);
mul_8x8bit m134 (image[72],filter[8],mul_out[44][2]);

adder_8bit ad14 (mul_out[42][0],mul_out[42][1],mul_out[42][2],mul_out[43][0],mul_out[43][1],mul_out[43][2],mul_out[44][0],mul_out[44][1],mul_out[44][2],conv_out[14]);



mul_8x8bit m135 (image[15],filter[0],mul_out[45][0]);
mul_8x8bit m136 (image[16],filter[1],mul_out[45][1]);
mul_8x8bit m137 (image[17],filter[2],mul_out[45][2]);
mul_8x8bit m138 (image[43],filter[3],mul_out[46][0]);
mul_8x8bit m139 (image[44],filter[4],mul_out[46][1]);
mul_8x8bit m140 (image[45],filter[5],mul_out[46][2]);
mul_8x8bit m141 (image[71],filter[6],mul_out[47][0]);
mul_8x8bit m142 (image[72],filter[7],mul_out[47][1]);
mul_8x8bit m143 (image[73],filter[8],mul_out[47][2]);

adder_8bit ad15 (mul_out[45][0],mul_out[45][1],mul_out[45][2],mul_out[46][0],mul_out[46][1],mul_out[46][2],mul_out[47][0],mul_out[47][1],mul_out[47][2],conv_out[15]);



mul_8x8bit m144 (image[16],filter[0],mul_out[48][0]);
mul_8x8bit m145 (image[17],filter[1],mul_out[48][1]);
mul_8x8bit m146 (image[18],filter[2],mul_out[48][2]);
mul_8x8bit m147 (image[44],filter[3],mul_out[49][0]);
mul_8x8bit m148 (image[45],filter[4],mul_out[49][1]);
mul_8x8bit m149 (image[46],filter[5],mul_out[49][2]);
mul_8x8bit m150 (image[72],filter[6],mul_out[50][0]);
mul_8x8bit m151 (image[73],filter[7],mul_out[50][1]);
mul_8x8bit m152 (image[74],filter[8],mul_out[50][2]);

adder_8bit ad16 (mul_out[48][0],mul_out[48][1],mul_out[48][2],mul_out[49][0],mul_out[49][1],mul_out[49][2],mul_out[50][0],mul_out[50][1],mul_out[50][2],conv_out[16]);



mul_8x8bit m153 (image[17],filter[0],mul_out[51][0]);
mul_8x8bit m154 (image[18],filter[1],mul_out[51][1]);
mul_8x8bit m155 (image[19],filter[2],mul_out[51][2]);
mul_8x8bit m156 (image[45],filter[3],mul_out[52][0]);
mul_8x8bit m157 (image[46],filter[4],mul_out[52][1]);
mul_8x8bit m158 (image[47],filter[5],mul_out[52][2]);
mul_8x8bit m159 (image[73],filter[6],mul_out[53][0]);
mul_8x8bit m160 (image[74],filter[7],mul_out[53][1]);
mul_8x8bit m161 (image[75],filter[8],mul_out[53][2]);

adder_8bit ad17 (mul_out[51][0],mul_out[51][1],mul_out[51][2],mul_out[52][0],mul_out[52][1],mul_out[52][2],mul_out[53][0],mul_out[53][1],mul_out[53][2],conv_out[17]);



mul_8x8bit m162 (image[18],filter[0],mul_out[54][0]);
mul_8x8bit m163 (image[19],filter[1],mul_out[54][1]);
mul_8x8bit m164 (image[20],filter[2],mul_out[54][2]);
mul_8x8bit m165 (image[46],filter[3],mul_out[55][0]);
mul_8x8bit m166 (image[47],filter[4],mul_out[55][1]);
mul_8x8bit m167 (image[48],filter[5],mul_out[55][2]);
mul_8x8bit m168 (image[74],filter[6],mul_out[56][0]);
mul_8x8bit m169 (image[75],filter[7],mul_out[56][1]);
mul_8x8bit m170 (image[76],filter[8],mul_out[56][2]);

adder_8bit ad18 (mul_out[54][0],mul_out[54][1],mul_out[54][2],mul_out[55][0],mul_out[55][1],mul_out[55][2],mul_out[56][0],mul_out[56][1],mul_out[56][2],conv_out[18]);



mul_8x8bit m171 (image[19],filter[0],mul_out[57][0]);
mul_8x8bit m172 (image[20],filter[1],mul_out[57][1]);
mul_8x8bit m173 (image[21],filter[2],mul_out[57][2]);
mul_8x8bit m174 (image[47],filter[3],mul_out[58][0]);
mul_8x8bit m175 (image[48],filter[4],mul_out[58][1]);
mul_8x8bit m176 (image[49],filter[5],mul_out[58][2]);
mul_8x8bit m177 (image[75],filter[6],mul_out[59][0]);
mul_8x8bit m178 (image[76],filter[7],mul_out[59][1]);
mul_8x8bit m179 (image[77],filter[8],mul_out[59][2]);

adder_8bit ad19 (mul_out[57][0],mul_out[57][1],mul_out[57][2],mul_out[58][0],mul_out[58][1],mul_out[58][2],mul_out[59][0],mul_out[59][1],mul_out[59][2],conv_out[19]);



mul_8x8bit m180 (image[20],filter[0],mul_out[60][0]);
mul_8x8bit m181 (image[21],filter[1],mul_out[60][1]);
mul_8x8bit m182 (image[22],filter[2],mul_out[60][2]);
mul_8x8bit m183 (image[48],filter[3],mul_out[61][0]);
mul_8x8bit m184 (image[49],filter[4],mul_out[61][1]);
mul_8x8bit m185 (image[50],filter[5],mul_out[61][2]);
mul_8x8bit m186 (image[76],filter[6],mul_out[62][0]);
mul_8x8bit m187 (image[77],filter[7],mul_out[62][1]);
mul_8x8bit m188 (image[78],filter[8],mul_out[62][2]);

adder_8bit ad20 (mul_out[60][0],mul_out[60][1],mul_out[60][2],mul_out[61][0],mul_out[61][1],mul_out[61][2],mul_out[62][0],mul_out[62][1],mul_out[62][2],conv_out[20]);



mul_8x8bit m189 (image[21],filter[0],mul_out[63][0]);
mul_8x8bit m190 (image[22],filter[1],mul_out[63][1]);
mul_8x8bit m191 (image[23],filter[2],mul_out[63][2]);
mul_8x8bit m192 (image[49],filter[3],mul_out[64][0]);
mul_8x8bit m193 (image[50],filter[4],mul_out[64][1]);
mul_8x8bit m194 (image[51],filter[5],mul_out[64][2]);
mul_8x8bit m195 (image[77],filter[6],mul_out[65][0]);
mul_8x8bit m196 (image[78],filter[7],mul_out[65][1]);
mul_8x8bit m197 (image[79],filter[8],mul_out[65][2]);

adder_8bit ad21 (mul_out[63][0],mul_out[63][1],mul_out[63][2],mul_out[64][0],mul_out[64][1],mul_out[64][2],mul_out[65][0],mul_out[65][1],mul_out[65][2],conv_out[21]);



mul_8x8bit m198 (image[22],filter[0],mul_out[66][0]);
mul_8x8bit m199 (image[23],filter[1],mul_out[66][1]);
mul_8x8bit m200 (image[24],filter[2],mul_out[66][2]);
mul_8x8bit m201 (image[50],filter[3],mul_out[67][0]);
mul_8x8bit m202 (image[51],filter[4],mul_out[67][1]);
mul_8x8bit m203 (image[52],filter[5],mul_out[67][2]);
mul_8x8bit m204 (image[78],filter[6],mul_out[68][0]);
mul_8x8bit m205 (image[79],filter[7],mul_out[68][1]);
mul_8x8bit m206 (image[80],filter[8],mul_out[68][2]);

adder_8bit ad22 (mul_out[66][0],mul_out[66][1],mul_out[66][2],mul_out[67][0],mul_out[67][1],mul_out[67][2],mul_out[68][0],mul_out[68][1],mul_out[68][2],conv_out[22]);



mul_8x8bit m207 (image[23],filter[0],mul_out[69][0]);
mul_8x8bit m208 (image[24],filter[1],mul_out[69][1]);
mul_8x8bit m209 (image[25],filter[2],mul_out[69][2]);
mul_8x8bit m210 (image[51],filter[3],mul_out[70][0]);
mul_8x8bit m211 (image[52],filter[4],mul_out[70][1]);
mul_8x8bit m212 (image[53],filter[5],mul_out[70][2]);
mul_8x8bit m213 (image[79],filter[6],mul_out[71][0]);
mul_8x8bit m214 (image[80],filter[7],mul_out[71][1]);
mul_8x8bit m215 (image[81],filter[8],mul_out[71][2]);

adder_8bit ad23 (mul_out[69][0],mul_out[69][1],mul_out[69][2],mul_out[70][0],mul_out[70][1],mul_out[70][2],mul_out[71][0],mul_out[71][1],mul_out[71][2],conv_out[23]);



mul_8x8bit m216 (image[24],filter[0],mul_out[72][0]);
mul_8x8bit m217 (image[25],filter[1],mul_out[72][1]);
mul_8x8bit m218 (image[26],filter[2],mul_out[72][2]);
mul_8x8bit m219 (image[52],filter[3],mul_out[73][0]);
mul_8x8bit m220 (image[53],filter[4],mul_out[73][1]);
mul_8x8bit m221 (image[54],filter[5],mul_out[73][2]);
mul_8x8bit m222 (image[80],filter[6],mul_out[74][0]);
mul_8x8bit m223 (image[81],filter[7],mul_out[74][1]);
mul_8x8bit m224 (image[82],filter[8],mul_out[74][2]);

adder_8bit ad24 (mul_out[72][0],mul_out[72][1],mul_out[72][2],mul_out[73][0],mul_out[73][1],mul_out[73][2],mul_out[74][0],mul_out[74][1],mul_out[74][2],conv_out[24]);



mul_8x8bit m225 (image[25],filter[0],mul_out[75][0]);
mul_8x8bit m226 (image[26],filter[1],mul_out[75][1]);
mul_8x8bit m227 (image[27],filter[2],mul_out[75][2]);
mul_8x8bit m228 (image[53],filter[3],mul_out[76][0]);
mul_8x8bit m229 (image[54],filter[4],mul_out[76][1]);
mul_8x8bit m230 (image[55],filter[5],mul_out[76][2]);
mul_8x8bit m231 (image[81],filter[6],mul_out[77][0]);
mul_8x8bit m232 (image[82],filter[7],mul_out[77][1]);
mul_8x8bit m233 (image[83],filter[8],mul_out[77][2]);

adder_8bit ad25 (mul_out[75][0],mul_out[75][1],mul_out[75][2],mul_out[76][0],mul_out[76][1],mul_out[76][2],mul_out[77][0],mul_out[77][1],mul_out[77][2],conv_out[25]);



mul_8x8bit m234 (image[28],filter[0],mul_out[78][1]);
mul_8x8bit m235 (image[29],filter[1],mul_out[78][2]);
mul_8x8bit m236 (image[30],filter[2],mul_out[78][3]);
mul_8x8bit m237 (image[56],filter[3],mul_out[79][1]);
mul_8x8bit m238 (image[57],filter[4],mul_out[79][2]);
mul_8x8bit m239 (image[58],filter[5],mul_out[79][3]);
mul_8x8bit m240 (image[84],filter[6],mul_out[80][1]);
mul_8x8bit m241 (image[85],filter[7],mul_out[80][2]);
mul_8x8bit m242 (image[86],filter[8],mul_out[80][3]);

adder_8bit ad26 (mul_out[78][1],mul_out[78][2],mul_out[78][3],mul_out[79][1],mul_out[79][2],mul_out[79][3],mul_out[80][1],mul_out[80][2],mul_out[80][3],conv_out[26]);



mul_8x8bit m243 (image[29],filter[0],mul_out[81][1]);
mul_8x8bit m244 (image[30],filter[1],mul_out[81][2]);
mul_8x8bit m245 (image[31],filter[2],mul_out[81][3]);
mul_8x8bit m246 (image[57],filter[3],mul_out[82][1]);
mul_8x8bit m247 (image[58],filter[4],mul_out[82][2]);
mul_8x8bit m248 (image[59],filter[5],mul_out[82][3]);
mul_8x8bit m249 (image[85],filter[6],mul_out[83][1]);
mul_8x8bit m250 (image[86],filter[7],mul_out[83][2]);
mul_8x8bit m251 (image[87],filter[8],mul_out[83][3]);

adder_8bit ad27 (mul_out[81][1],mul_out[81][2],mul_out[81][3],mul_out[82][1],mul_out[82][2],mul_out[82][3],mul_out[83][1],mul_out[83][2],mul_out[83][3],conv_out[27]);



mul_8x8bit m252 (image[30],filter[0],mul_out[84][1]);
mul_8x8bit m253 (image[31],filter[1],mul_out[84][2]);
mul_8x8bit m254 (image[32],filter[2],mul_out[84][3]);
mul_8x8bit m255 (image[58],filter[3],mul_out[85][1]);
mul_8x8bit m256 (image[59],filter[4],mul_out[85][2]);
mul_8x8bit m257 (image[60],filter[5],mul_out[85][3]);
mul_8x8bit m258 (image[86],filter[6],mul_out[86][1]);
mul_8x8bit m259 (image[87],filter[7],mul_out[86][2]);
mul_8x8bit m260 (image[88],filter[8],mul_out[86][3]);

adder_8bit ad28 (mul_out[84][1],mul_out[84][2],mul_out[84][3],mul_out[85][1],mul_out[85][2],mul_out[85][3],mul_out[86][1],mul_out[86][2],mul_out[86][3],conv_out[28]);



mul_8x8bit m261 (image[31],filter[0],mul_out[87][1]);
mul_8x8bit m262 (image[32],filter[1],mul_out[87][2]);
mul_8x8bit m263 (image[33],filter[2],mul_out[87][3]);
mul_8x8bit m264 (image[59],filter[3],mul_out[88][1]);
mul_8x8bit m265 (image[60],filter[4],mul_out[88][2]);
mul_8x8bit m266 (image[61],filter[5],mul_out[88][3]);
mul_8x8bit m267 (image[87],filter[6],mul_out[89][1]);
mul_8x8bit m268 (image[88],filter[7],mul_out[89][2]);
mul_8x8bit m269 (image[89],filter[8],mul_out[89][3]);

adder_8bit ad29 (mul_out[87][1],mul_out[87][2],mul_out[87][3],mul_out[88][1],mul_out[88][2],mul_out[88][3],mul_out[89][1],mul_out[89][2],mul_out[89][3],conv_out[29]);



mul_8x8bit m270 (image[32],filter[0],mul_out[90][1]);
mul_8x8bit m271 (image[33],filter[1],mul_out[90][2]);
mul_8x8bit m272 (image[34],filter[2],mul_out[90][3]);
mul_8x8bit m273 (image[60],filter[3],mul_out[91][1]);
mul_8x8bit m274 (image[61],filter[4],mul_out[91][2]);
mul_8x8bit m275 (image[62],filter[5],mul_out[91][3]);
mul_8x8bit m276 (image[88],filter[6],mul_out[92][1]);
mul_8x8bit m277 (image[89],filter[7],mul_out[92][2]);
mul_8x8bit m278 (image[90],filter[8],mul_out[92][3]);

adder_8bit ad30 (mul_out[90][1],mul_out[90][2],mul_out[90][3],mul_out[91][1],mul_out[91][2],mul_out[91][3],mul_out[92][1],mul_out[92][2],mul_out[92][3],conv_out[30]);



mul_8x8bit m279 (image[33],filter[0],mul_out[93][1]);
mul_8x8bit m280 (image[34],filter[1],mul_out[93][2]);
mul_8x8bit m281 (image[35],filter[2],mul_out[93][3]);
mul_8x8bit m282 (image[61],filter[3],mul_out[94][1]);
mul_8x8bit m283 (image[62],filter[4],mul_out[94][2]);
mul_8x8bit m284 (image[63],filter[5],mul_out[94][3]);
mul_8x8bit m285 (image[89],filter[6],mul_out[95][1]);
mul_8x8bit m286 (image[90],filter[7],mul_out[95][2]);
mul_8x8bit m287 (image[91],filter[8],mul_out[95][3]);

adder_8bit ad31 (mul_out[93][1],mul_out[93][2],mul_out[93][3],mul_out[94][1],mul_out[94][2],mul_out[94][3],mul_out[95][1],mul_out[95][2],mul_out[95][3],conv_out[31]);



mul_8x8bit m288 (image[34],filter[0],mul_out[96][1]);
mul_8x8bit m289 (image[35],filter[1],mul_out[96][2]);
mul_8x8bit m290 (image[36],filter[2],mul_out[96][3]);
mul_8x8bit m291 (image[62],filter[3],mul_out[97][1]);
mul_8x8bit m292 (image[63],filter[4],mul_out[97][2]);
mul_8x8bit m293 (image[64],filter[5],mul_out[97][3]);
mul_8x8bit m294 (image[90],filter[6],mul_out[98][1]);
mul_8x8bit m295 (image[91],filter[7],mul_out[98][2]);
mul_8x8bit m296 (image[92],filter[8],mul_out[98][3]);

adder_8bit ad32 (mul_out[96][1],mul_out[96][2],mul_out[96][3],mul_out[97][1],mul_out[97][2],mul_out[97][3],mul_out[98][1],mul_out[98][2],mul_out[98][3],conv_out[32]);



mul_8x8bit m297 (image[35],filter[0],mul_out[99][1]);
mul_8x8bit m298 (image[36],filter[1],mul_out[99][2]);
mul_8x8bit m299 (image[37],filter[2],mul_out[99][3]);
mul_8x8bit m300 (image[63],filter[3],mul_out[100][1]);
mul_8x8bit m301 (image[64],filter[4],mul_out[100][2]);
mul_8x8bit m302 (image[65],filter[5],mul_out[100][3]);
mul_8x8bit m303 (image[91],filter[6],mul_out[101][1]);
mul_8x8bit m304 (image[92],filter[7],mul_out[101][2]);
mul_8x8bit m305 (image[93],filter[8],mul_out[101][3]);

adder_8bit ad33 (mul_out[99][1],mul_out[99][2],mul_out[99][3],mul_out[100][1],mul_out[100][2],mul_out[100][3],mul_out[101][1],mul_out[101][2],mul_out[101][3],conv_out[33]);



mul_8x8bit m306 (image[36],filter[0],mul_out[102][1]);
mul_8x8bit m307 (image[37],filter[1],mul_out[102][2]);
mul_8x8bit m308 (image[38],filter[2],mul_out[102][3]);
mul_8x8bit m309 (image[64],filter[3],mul_out[103][1]);
mul_8x8bit m310 (image[65],filter[4],mul_out[103][2]);
mul_8x8bit m311 (image[66],filter[5],mul_out[103][3]);
mul_8x8bit m312 (image[92],filter[6],mul_out[104][1]);
mul_8x8bit m313 (image[93],filter[7],mul_out[104][2]);
mul_8x8bit m314 (image[94],filter[8],mul_out[104][3]);

adder_8bit ad34 (mul_out[102][1],mul_out[102][2],mul_out[102][3],mul_out[103][1],mul_out[103][2],mul_out[103][3],mul_out[104][1],mul_out[104][2],mul_out[104][3],conv_out[34]);



mul_8x8bit m315 (image[37],filter[0],mul_out[105][1]);
mul_8x8bit m316 (image[38],filter[1],mul_out[105][2]);
mul_8x8bit m317 (image[39],filter[2],mul_out[105][3]);
mul_8x8bit m318 (image[65],filter[3],mul_out[106][1]);
mul_8x8bit m319 (image[66],filter[4],mul_out[106][2]);
mul_8x8bit m320 (image[67],filter[5],mul_out[106][3]);
mul_8x8bit m321 (image[93],filter[6],mul_out[107][1]);
mul_8x8bit m322 (image[94],filter[7],mul_out[107][2]);
mul_8x8bit m323 (image[95],filter[8],mul_out[107][3]);

adder_8bit ad35 (mul_out[105][1],mul_out[105][2],mul_out[105][3],mul_out[106][1],mul_out[106][2],mul_out[106][3],mul_out[107][1],mul_out[107][2],mul_out[107][3],conv_out[35]);



mul_8x8bit m324 (image[38],filter[0],mul_out[108][1]);
mul_8x8bit m325 (image[39],filter[1],mul_out[108][2]);
mul_8x8bit m326 (image[40],filter[2],mul_out[108][3]);
mul_8x8bit m327 (image[66],filter[3],mul_out[109][1]);
mul_8x8bit m328 (image[67],filter[4],mul_out[109][2]);
mul_8x8bit m329 (image[68],filter[5],mul_out[109][3]);
mul_8x8bit m330 (image[94],filter[6],mul_out[110][1]);
mul_8x8bit m331 (image[95],filter[7],mul_out[110][2]);
mul_8x8bit m332 (image[96],filter[8],mul_out[110][3]);

adder_8bit ad36 (mul_out[108][1],mul_out[108][2],mul_out[108][3],mul_out[109][1],mul_out[109][2],mul_out[109][3],mul_out[110][1],mul_out[110][2],mul_out[110][3],conv_out[36]);



mul_8x8bit m333 (image[39],filter[0],mul_out[111][1]);
mul_8x8bit m334 (image[40],filter[1],mul_out[111][2]);
mul_8x8bit m335 (image[41],filter[2],mul_out[111][3]);
mul_8x8bit m336 (image[67],filter[3],mul_out[112][1]);
mul_8x8bit m337 (image[68],filter[4],mul_out[112][2]);
mul_8x8bit m338 (image[69],filter[5],mul_out[112][3]);
mul_8x8bit m339 (image[95],filter[6],mul_out[113][1]);
mul_8x8bit m340 (image[96],filter[7],mul_out[113][2]);
mul_8x8bit m341 (image[97],filter[8],mul_out[113][3]);

adder_8bit ad37 (mul_out[111][1],mul_out[111][2],mul_out[111][3],mul_out[112][1],mul_out[112][2],mul_out[112][3],mul_out[113][1],mul_out[113][2],mul_out[113][3],conv_out[37]);



mul_8x8bit m342 (image[40],filter[0],mul_out[114][1]);
mul_8x8bit m343 (image[41],filter[1],mul_out[114][2]);
mul_8x8bit m344 (image[42],filter[2],mul_out[114][3]);
mul_8x8bit m345 (image[68],filter[3],mul_out[115][1]);
mul_8x8bit m346 (image[69],filter[4],mul_out[115][2]);
mul_8x8bit m347 (image[70],filter[5],mul_out[115][3]);
mul_8x8bit m348 (image[96],filter[6],mul_out[116][1]);
mul_8x8bit m349 (image[97],filter[7],mul_out[116][2]);
mul_8x8bit m350 (image[98],filter[8],mul_out[116][3]);

adder_8bit ad38 (mul_out[114][1],mul_out[114][2],mul_out[114][3],mul_out[115][1],mul_out[115][2],mul_out[115][3],mul_out[116][1],mul_out[116][2],mul_out[116][3],conv_out[38]);



mul_8x8bit m351 (image[41],filter[0],mul_out[117][1]);
mul_8x8bit m352 (image[42],filter[1],mul_out[117][2]);
mul_8x8bit m353 (image[43],filter[2],mul_out[117][3]);
mul_8x8bit m354 (image[69],filter[3],mul_out[118][1]);
mul_8x8bit m355 (image[70],filter[4],mul_out[118][2]);
mul_8x8bit m356 (image[71],filter[5],mul_out[118][3]);
mul_8x8bit m357 (image[97],filter[6],mul_out[119][1]);
mul_8x8bit m358 (image[98],filter[7],mul_out[119][2]);
mul_8x8bit m359 (image[99],filter[8],mul_out[119][3]);

adder_8bit ad39 (mul_out[117][1],mul_out[117][2],mul_out[117][3],mul_out[118][1],mul_out[118][2],mul_out[118][3],mul_out[119][1],mul_out[119][2],mul_out[119][3],conv_out[39]);



mul_8x8bit m360 (image[42],filter[0],mul_out[120][1]);
mul_8x8bit m361 (image[43],filter[1],mul_out[120][2]);
mul_8x8bit m362 (image[44],filter[2],mul_out[120][3]);
mul_8x8bit m363 (image[70],filter[3],mul_out[121][1]);
mul_8x8bit m364 (image[71],filter[4],mul_out[121][2]);
mul_8x8bit m365 (image[72],filter[5],mul_out[121][3]);
mul_8x8bit m366 (image[98],filter[6],mul_out[122][1]);
mul_8x8bit m367 (image[99],filter[7],mul_out[122][2]);
mul_8x8bit m368 (image[100],filter[8],mul_out[122][3]);

adder_8bit ad40 (mul_out[120][1],mul_out[120][2],mul_out[120][3],mul_out[121][1],mul_out[121][2],mul_out[121][3],mul_out[122][1],mul_out[122][2],mul_out[122][3],conv_out[40]);



mul_8x8bit m369 (image[43],filter[0],mul_out[123][1]);
mul_8x8bit m370 (image[44],filter[1],mul_out[123][2]);
mul_8x8bit m371 (image[45],filter[2],mul_out[123][3]);
mul_8x8bit m372 (image[71],filter[3],mul_out[124][1]);
mul_8x8bit m373 (image[72],filter[4],mul_out[124][2]);
mul_8x8bit m374 (image[73],filter[5],mul_out[124][3]);
mul_8x8bit m375 (image[99],filter[6],mul_out[125][1]);
mul_8x8bit m376 (image[100],filter[7],mul_out[125][2]);
mul_8x8bit m377 (image[101],filter[8],mul_out[125][3]);

adder_8bit ad41 (mul_out[123][1],mul_out[123][2],mul_out[123][3],mul_out[124][1],mul_out[124][2],mul_out[124][3],mul_out[125][1],mul_out[125][2],mul_out[125][3],conv_out[41]);



mul_8x8bit m378 (image[44],filter[0],mul_out[126][1]);
mul_8x8bit m379 (image[45],filter[1],mul_out[126][2]);
mul_8x8bit m380 (image[46],filter[2],mul_out[126][3]);
mul_8x8bit m381 (image[72],filter[3],mul_out[127][1]);
mul_8x8bit m382 (image[73],filter[4],mul_out[127][2]);
mul_8x8bit m383 (image[74],filter[5],mul_out[127][3]);
mul_8x8bit m384 (image[100],filter[6],mul_out[128][1]);
mul_8x8bit m385 (image[101],filter[7],mul_out[128][2]);
mul_8x8bit m386 (image[102],filter[8],mul_out[128][3]);

adder_8bit ad42 (mul_out[126][1],mul_out[126][2],mul_out[126][3],mul_out[127][1],mul_out[127][2],mul_out[127][3],mul_out[128][1],mul_out[128][2],mul_out[128][3],conv_out[42]);



mul_8x8bit m387 (image[45],filter[0],mul_out[129][1]);
mul_8x8bit m388 (image[46],filter[1],mul_out[129][2]);
mul_8x8bit m389 (image[47],filter[2],mul_out[129][3]);
mul_8x8bit m390 (image[73],filter[3],mul_out[130][1]);
mul_8x8bit m391 (image[74],filter[4],mul_out[130][2]);
mul_8x8bit m392 (image[75],filter[5],mul_out[130][3]);
mul_8x8bit m393 (image[101],filter[6],mul_out[131][1]);
mul_8x8bit m394 (image[102],filter[7],mul_out[131][2]);
mul_8x8bit m395 (image[103],filter[8],mul_out[131][3]);

adder_8bit ad43 (mul_out[129][1],mul_out[129][2],mul_out[129][3],mul_out[130][1],mul_out[130][2],mul_out[130][3],mul_out[131][1],mul_out[131][2],mul_out[131][3],conv_out[43]);



mul_8x8bit m396 (image[46],filter[0],mul_out[132][1]);
mul_8x8bit m397 (image[47],filter[1],mul_out[132][2]);
mul_8x8bit m398 (image[48],filter[2],mul_out[132][3]);
mul_8x8bit m399 (image[74],filter[3],mul_out[133][1]);
mul_8x8bit m400 (image[75],filter[4],mul_out[133][2]);
mul_8x8bit m401 (image[76],filter[5],mul_out[133][3]);
mul_8x8bit m402 (image[102],filter[6],mul_out[134][1]);
mul_8x8bit m403 (image[103],filter[7],mul_out[134][2]);
mul_8x8bit m404 (image[104],filter[8],mul_out[134][3]);

adder_8bit ad44 (mul_out[132][1],mul_out[132][2],mul_out[132][3],mul_out[133][1],mul_out[133][2],mul_out[133][3],mul_out[134][1],mul_out[134][2],mul_out[134][3],conv_out[44]);



mul_8x8bit m405 (image[47],filter[0],mul_out[135][1]);
mul_8x8bit m406 (image[48],filter[1],mul_out[135][2]);
mul_8x8bit m407 (image[49],filter[2],mul_out[135][3]);
mul_8x8bit m408 (image[75],filter[3],mul_out[136][1]);
mul_8x8bit m409 (image[76],filter[4],mul_out[136][2]);
mul_8x8bit m410 (image[77],filter[5],mul_out[136][3]);
mul_8x8bit m411 (image[103],filter[6],mul_out[137][1]);
mul_8x8bit m412 (image[104],filter[7],mul_out[137][2]);
mul_8x8bit m413 (image[105],filter[8],mul_out[137][3]);

adder_8bit ad45 (mul_out[135][1],mul_out[135][2],mul_out[135][3],mul_out[136][1],mul_out[136][2],mul_out[136][3],mul_out[137][1],mul_out[137][2],mul_out[137][3],conv_out[45]);



mul_8x8bit m414 (image[48],filter[0],mul_out[138][1]);
mul_8x8bit m415 (image[49],filter[1],mul_out[138][2]);
mul_8x8bit m416 (image[50],filter[2],mul_out[138][3]);
mul_8x8bit m417 (image[76],filter[3],mul_out[139][1]);
mul_8x8bit m418 (image[77],filter[4],mul_out[139][2]);
mul_8x8bit m419 (image[78],filter[5],mul_out[139][3]);
mul_8x8bit m420 (image[104],filter[6],mul_out[140][1]);
mul_8x8bit m421 (image[105],filter[7],mul_out[140][2]);
mul_8x8bit m422 (image[106],filter[8],mul_out[140][3]);

adder_8bit ad46 (mul_out[138][1],mul_out[138][2],mul_out[138][3],mul_out[139][1],mul_out[139][2],mul_out[139][3],mul_out[140][1],mul_out[140][2],mul_out[140][3],conv_out[46]);



mul_8x8bit m423 (image[49],filter[0],mul_out[141][1]);
mul_8x8bit m424 (image[50],filter[1],mul_out[141][2]);
mul_8x8bit m425 (image[51],filter[2],mul_out[141][3]);
mul_8x8bit m426 (image[77],filter[3],mul_out[142][1]);
mul_8x8bit m427 (image[78],filter[4],mul_out[142][2]);
mul_8x8bit m428 (image[79],filter[5],mul_out[142][3]);
mul_8x8bit m429 (image[105],filter[6],mul_out[143][1]);
mul_8x8bit m430 (image[106],filter[7],mul_out[143][2]);
mul_8x8bit m431 (image[107],filter[8],mul_out[143][3]);

adder_8bit ad47 (mul_out[141][1],mul_out[141][2],mul_out[141][3],mul_out[142][1],mul_out[142][2],mul_out[142][3],mul_out[143][1],mul_out[143][2],mul_out[143][3],conv_out[47]);



mul_8x8bit m432 (image[50],filter[0],mul_out[144][1]);
mul_8x8bit m433 (image[51],filter[1],mul_out[144][2]);
mul_8x8bit m434 (image[52],filter[2],mul_out[144][3]);
mul_8x8bit m435 (image[78],filter[3],mul_out[145][1]);
mul_8x8bit m436 (image[79],filter[4],mul_out[145][2]);
mul_8x8bit m437 (image[80],filter[5],mul_out[145][3]);
mul_8x8bit m438 (image[106],filter[6],mul_out[146][1]);
mul_8x8bit m439 (image[107],filter[7],mul_out[146][2]);
mul_8x8bit m440 (image[108],filter[8],mul_out[146][3]);

adder_8bit ad48 (mul_out[144][1],mul_out[144][2],mul_out[144][3],mul_out[145][1],mul_out[145][2],mul_out[145][3],mul_out[146][1],mul_out[146][2],mul_out[146][3],conv_out[48]);



mul_8x8bit m441 (image[51],filter[0],mul_out[147][1]);
mul_8x8bit m442 (image[52],filter[1],mul_out[147][2]);
mul_8x8bit m443 (image[53],filter[2],mul_out[147][3]);
mul_8x8bit m444 (image[79],filter[3],mul_out[148][1]);
mul_8x8bit m445 (image[80],filter[4],mul_out[148][2]);
mul_8x8bit m446 (image[81],filter[5],mul_out[148][3]);
mul_8x8bit m447 (image[107],filter[6],mul_out[149][1]);
mul_8x8bit m448 (image[108],filter[7],mul_out[149][2]);
mul_8x8bit m449 (image[109],filter[8],mul_out[149][3]);

adder_8bit ad49 (mul_out[147][1],mul_out[147][2],mul_out[147][3],mul_out[148][1],mul_out[148][2],mul_out[148][3],mul_out[149][1],mul_out[149][2],mul_out[149][3],conv_out[49]);



mul_8x8bit m450 (image[52],filter[0],mul_out[150][1]);
mul_8x8bit m451 (image[53],filter[1],mul_out[150][2]);
mul_8x8bit m452 (image[54],filter[2],mul_out[150][3]);
mul_8x8bit m453 (image[80],filter[3],mul_out[151][1]);
mul_8x8bit m454 (image[81],filter[4],mul_out[151][2]);
mul_8x8bit m455 (image[82],filter[5],mul_out[151][3]);
mul_8x8bit m456 (image[108],filter[6],mul_out[152][1]);
mul_8x8bit m457 (image[109],filter[7],mul_out[152][2]);
mul_8x8bit m458 (image[110],filter[8],mul_out[152][3]);

adder_8bit ad50 (mul_out[150][1],mul_out[150][2],mul_out[150][3],mul_out[151][1],mul_out[151][2],mul_out[151][3],mul_out[152][1],mul_out[152][2],mul_out[152][3],conv_out[50]);



mul_8x8bit m459 (image[53],filter[0],mul_out[153][1]);
mul_8x8bit m460 (image[54],filter[1],mul_out[153][2]);
mul_8x8bit m461 (image[55],filter[2],mul_out[153][3]);
mul_8x8bit m462 (image[81],filter[3],mul_out[154][1]);
mul_8x8bit m463 (image[82],filter[4],mul_out[154][2]);
mul_8x8bit m464 (image[83],filter[5],mul_out[154][3]);
mul_8x8bit m465 (image[109],filter[6],mul_out[155][1]);
mul_8x8bit m466 (image[110],filter[7],mul_out[155][2]);
mul_8x8bit m467 (image[111],filter[8],mul_out[155][3]);

adder_8bit ad51 (mul_out[153][1],mul_out[153][2],mul_out[153][3],mul_out[154][1],mul_out[154][2],mul_out[154][3],mul_out[155][1],mul_out[155][2],mul_out[155][3],conv_out[51]);



mul_8x8bit m468 (image[56],filter[0],mul_out[156][2]);
mul_8x8bit m469 (image[57],filter[1],mul_out[156][3]);
mul_8x8bit m470 (image[58],filter[2],mul_out[156][4]);
mul_8x8bit m471 (image[84],filter[3],mul_out[157][2]);
mul_8x8bit m472 (image[85],filter[4],mul_out[157][3]);
mul_8x8bit m473 (image[86],filter[5],mul_out[157][4]);
mul_8x8bit m474 (image[112],filter[6],mul_out[158][2]);
mul_8x8bit m475 (image[113],filter[7],mul_out[158][3]);
mul_8x8bit m476 (image[114],filter[8],mul_out[158][4]);

adder_8bit ad52 (mul_out[156][2],mul_out[156][3],mul_out[156][4],mul_out[157][2],mul_out[157][3],mul_out[157][4],mul_out[158][2],mul_out[158][3],mul_out[158][4],conv_out[52]);



mul_8x8bit m477 (image[57],filter[0],mul_out[159][2]);
mul_8x8bit m478 (image[58],filter[1],mul_out[159][3]);
mul_8x8bit m479 (image[59],filter[2],mul_out[159][4]);
mul_8x8bit m480 (image[85],filter[3],mul_out[160][2]);
mul_8x8bit m481 (image[86],filter[4],mul_out[160][3]);
mul_8x8bit m482 (image[87],filter[5],mul_out[160][4]);
mul_8x8bit m483 (image[113],filter[6],mul_out[161][2]);
mul_8x8bit m484 (image[114],filter[7],mul_out[161][3]);
mul_8x8bit m485 (image[115],filter[8],mul_out[161][4]);

adder_8bit ad53 (mul_out[159][2],mul_out[159][3],mul_out[159][4],mul_out[160][2],mul_out[160][3],mul_out[160][4],mul_out[161][2],mul_out[161][3],mul_out[161][4],conv_out[53]);



mul_8x8bit m486 (image[58],filter[0],mul_out[162][2]);
mul_8x8bit m487 (image[59],filter[1],mul_out[162][3]);
mul_8x8bit m488 (image[60],filter[2],mul_out[162][4]);
mul_8x8bit m489 (image[86],filter[3],mul_out[163][2]);
mul_8x8bit m490 (image[87],filter[4],mul_out[163][3]);
mul_8x8bit m491 (image[88],filter[5],mul_out[163][4]);
mul_8x8bit m492 (image[114],filter[6],mul_out[164][2]);
mul_8x8bit m493 (image[115],filter[7],mul_out[164][3]);
mul_8x8bit m494 (image[116],filter[8],mul_out[164][4]);

adder_8bit ad54 (mul_out[162][2],mul_out[162][3],mul_out[162][4],mul_out[163][2],mul_out[163][3],mul_out[163][4],mul_out[164][2],mul_out[164][3],mul_out[164][4],conv_out[54]);



mul_8x8bit m495 (image[59],filter[0],mul_out[165][2]);
mul_8x8bit m496 (image[60],filter[1],mul_out[165][3]);
mul_8x8bit m497 (image[61],filter[2],mul_out[165][4]);
mul_8x8bit m498 (image[87],filter[3],mul_out[166][2]);
mul_8x8bit m499 (image[88],filter[4],mul_out[166][3]);
mul_8x8bit m500 (image[89],filter[5],mul_out[166][4]);
mul_8x8bit m501 (image[115],filter[6],mul_out[167][2]);
mul_8x8bit m502 (image[116],filter[7],mul_out[167][3]);
mul_8x8bit m503 (image[117],filter[8],mul_out[167][4]);

adder_8bit ad55 (mul_out[165][2],mul_out[165][3],mul_out[165][4],mul_out[166][2],mul_out[166][3],mul_out[166][4],mul_out[167][2],mul_out[167][3],mul_out[167][4],conv_out[55]);



mul_8x8bit m504 (image[60],filter[0],mul_out[168][2]);
mul_8x8bit m505 (image[61],filter[1],mul_out[168][3]);
mul_8x8bit m506 (image[62],filter[2],mul_out[168][4]);
mul_8x8bit m507 (image[88],filter[3],mul_out[169][2]);
mul_8x8bit m508 (image[89],filter[4],mul_out[169][3]);
mul_8x8bit m509 (image[90],filter[5],mul_out[169][4]);
mul_8x8bit m510 (image[116],filter[6],mul_out[170][2]);
mul_8x8bit m511 (image[117],filter[7],mul_out[170][3]);
mul_8x8bit m512 (image[118],filter[8],mul_out[170][4]);

adder_8bit ad56 (mul_out[168][2],mul_out[168][3],mul_out[168][4],mul_out[169][2],mul_out[169][3],mul_out[169][4],mul_out[170][2],mul_out[170][3],mul_out[170][4],conv_out[56]);



mul_8x8bit m513 (image[61],filter[0],mul_out[171][2]);
mul_8x8bit m514 (image[62],filter[1],mul_out[171][3]);
mul_8x8bit m515 (image[63],filter[2],mul_out[171][4]);
mul_8x8bit m516 (image[89],filter[3],mul_out[172][2]);
mul_8x8bit m517 (image[90],filter[4],mul_out[172][3]);
mul_8x8bit m518 (image[91],filter[5],mul_out[172][4]);
mul_8x8bit m519 (image[117],filter[6],mul_out[173][2]);
mul_8x8bit m520 (image[118],filter[7],mul_out[173][3]);
mul_8x8bit m521 (image[119],filter[8],mul_out[173][4]);

adder_8bit ad57 (mul_out[171][2],mul_out[171][3],mul_out[171][4],mul_out[172][2],mul_out[172][3],mul_out[172][4],mul_out[173][2],mul_out[173][3],mul_out[173][4],conv_out[57]);



mul_8x8bit m522 (image[62],filter[0],mul_out[174][2]);
mul_8x8bit m523 (image[63],filter[1],mul_out[174][3]);
mul_8x8bit m524 (image[64],filter[2],mul_out[174][4]);
mul_8x8bit m525 (image[90],filter[3],mul_out[175][2]);
mul_8x8bit m526 (image[91],filter[4],mul_out[175][3]);
mul_8x8bit m527 (image[92],filter[5],mul_out[175][4]);
mul_8x8bit m528 (image[118],filter[6],mul_out[176][2]);
mul_8x8bit m529 (image[119],filter[7],mul_out[176][3]);
mul_8x8bit m530 (image[120],filter[8],mul_out[176][4]);

adder_8bit ad58 (mul_out[174][2],mul_out[174][3],mul_out[174][4],mul_out[175][2],mul_out[175][3],mul_out[175][4],mul_out[176][2],mul_out[176][3],mul_out[176][4],conv_out[58]);



mul_8x8bit m531 (image[63],filter[0],mul_out[177][2]);
mul_8x8bit m532 (image[64],filter[1],mul_out[177][3]);
mul_8x8bit m533 (image[65],filter[2],mul_out[177][4]);
mul_8x8bit m534 (image[91],filter[3],mul_out[178][2]);
mul_8x8bit m535 (image[92],filter[4],mul_out[178][3]);
mul_8x8bit m536 (image[93],filter[5],mul_out[178][4]);
mul_8x8bit m537 (image[119],filter[6],mul_out[179][2]);
mul_8x8bit m538 (image[120],filter[7],mul_out[179][3]);
mul_8x8bit m539 (image[121],filter[8],mul_out[179][4]);

adder_8bit ad59 (mul_out[177][2],mul_out[177][3],mul_out[177][4],mul_out[178][2],mul_out[178][3],mul_out[178][4],mul_out[179][2],mul_out[179][3],mul_out[179][4],conv_out[59]);



mul_8x8bit m540 (image[64],filter[0],mul_out[180][2]);
mul_8x8bit m541 (image[65],filter[1],mul_out[180][3]);
mul_8x8bit m542 (image[66],filter[2],mul_out[180][4]);
mul_8x8bit m543 (image[92],filter[3],mul_out[181][2]);
mul_8x8bit m544 (image[93],filter[4],mul_out[181][3]);
mul_8x8bit m545 (image[94],filter[5],mul_out[181][4]);
mul_8x8bit m546 (image[120],filter[6],mul_out[182][2]);
mul_8x8bit m547 (image[121],filter[7],mul_out[182][3]);
mul_8x8bit m548 (image[122],filter[8],mul_out[182][4]);

adder_8bit ad60 (mul_out[180][2],mul_out[180][3],mul_out[180][4],mul_out[181][2],mul_out[181][3],mul_out[181][4],mul_out[182][2],mul_out[182][3],mul_out[182][4],conv_out[60]);



mul_8x8bit m549 (image[65],filter[0],mul_out[183][2]);
mul_8x8bit m550 (image[66],filter[1],mul_out[183][3]);
mul_8x8bit m551 (image[67],filter[2],mul_out[183][4]);
mul_8x8bit m552 (image[93],filter[3],mul_out[184][2]);
mul_8x8bit m553 (image[94],filter[4],mul_out[184][3]);
mul_8x8bit m554 (image[95],filter[5],mul_out[184][4]);
mul_8x8bit m555 (image[121],filter[6],mul_out[185][2]);
mul_8x8bit m556 (image[122],filter[7],mul_out[185][3]);
mul_8x8bit m557 (image[123],filter[8],mul_out[185][4]);

adder_8bit ad61 (mul_out[183][2],mul_out[183][3],mul_out[183][4],mul_out[184][2],mul_out[184][3],mul_out[184][4],mul_out[185][2],mul_out[185][3],mul_out[185][4],conv_out[61]);



mul_8x8bit m558 (image[66],filter[0],mul_out[186][2]);
mul_8x8bit m559 (image[67],filter[1],mul_out[186][3]);
mul_8x8bit m560 (image[68],filter[2],mul_out[186][4]);
mul_8x8bit m561 (image[94],filter[3],mul_out[187][2]);
mul_8x8bit m562 (image[95],filter[4],mul_out[187][3]);
mul_8x8bit m563 (image[96],filter[5],mul_out[187][4]);
mul_8x8bit m564 (image[122],filter[6],mul_out[188][2]);
mul_8x8bit m565 (image[123],filter[7],mul_out[188][3]);
mul_8x8bit m566 (image[124],filter[8],mul_out[188][4]);

adder_8bit ad62 (mul_out[186][2],mul_out[186][3],mul_out[186][4],mul_out[187][2],mul_out[187][3],mul_out[187][4],mul_out[188][2],mul_out[188][3],mul_out[188][4],conv_out[62]);



mul_8x8bit m567 (image[67],filter[0],mul_out[189][2]);
mul_8x8bit m568 (image[68],filter[1],mul_out[189][3]);
mul_8x8bit m569 (image[69],filter[2],mul_out[189][4]);
mul_8x8bit m570 (image[95],filter[3],mul_out[190][2]);
mul_8x8bit m571 (image[96],filter[4],mul_out[190][3]);
mul_8x8bit m572 (image[97],filter[5],mul_out[190][4]);
mul_8x8bit m573 (image[123],filter[6],mul_out[191][2]);
mul_8x8bit m574 (image[124],filter[7],mul_out[191][3]);
mul_8x8bit m575 (image[125],filter[8],mul_out[191][4]);

adder_8bit ad63 (mul_out[189][2],mul_out[189][3],mul_out[189][4],mul_out[190][2],mul_out[190][3],mul_out[190][4],mul_out[191][2],mul_out[191][3],mul_out[191][4],conv_out[63]);



mul_8x8bit m576 (image[68],filter[0],mul_out[192][2]);
mul_8x8bit m577 (image[69],filter[1],mul_out[192][3]);
mul_8x8bit m578 (image[70],filter[2],mul_out[192][4]);
mul_8x8bit m579 (image[96],filter[3],mul_out[193][2]);
mul_8x8bit m580 (image[97],filter[4],mul_out[193][3]);
mul_8x8bit m581 (image[98],filter[5],mul_out[193][4]);
mul_8x8bit m582 (image[124],filter[6],mul_out[194][2]);
mul_8x8bit m583 (image[125],filter[7],mul_out[194][3]);
mul_8x8bit m584 (image[126],filter[8],mul_out[194][4]);

adder_8bit ad64 (mul_out[192][2],mul_out[192][3],mul_out[192][4],mul_out[193][2],mul_out[193][3],mul_out[193][4],mul_out[194][2],mul_out[194][3],mul_out[194][4],conv_out[64]);



mul_8x8bit m585 (image[69],filter[0],mul_out[195][2]);
mul_8x8bit m586 (image[70],filter[1],mul_out[195][3]);
mul_8x8bit m587 (image[71],filter[2],mul_out[195][4]);
mul_8x8bit m588 (image[97],filter[3],mul_out[196][2]);
mul_8x8bit m589 (image[98],filter[4],mul_out[196][3]);
mul_8x8bit m590 (image[99],filter[5],mul_out[196][4]);
mul_8x8bit m591 (image[125],filter[6],mul_out[197][2]);
mul_8x8bit m592 (image[126],filter[7],mul_out[197][3]);
mul_8x8bit m593 (image[127],filter[8],mul_out[197][4]);

adder_8bit ad65 (mul_out[195][2],mul_out[195][3],mul_out[195][4],mul_out[196][2],mul_out[196][3],mul_out[196][4],mul_out[197][2],mul_out[197][3],mul_out[197][4],conv_out[65]);



mul_8x8bit m594 (image[70],filter[0],mul_out[198][2]);
mul_8x8bit m595 (image[71],filter[1],mul_out[198][3]);
mul_8x8bit m596 (image[72],filter[2],mul_out[198][4]);
mul_8x8bit m597 (image[98],filter[3],mul_out[199][2]);
mul_8x8bit m598 (image[99],filter[4],mul_out[199][3]);
mul_8x8bit m599 (image[100],filter[5],mul_out[199][4]);
mul_8x8bit m600 (image[126],filter[6],mul_out[200][2]);
mul_8x8bit m601 (image[127],filter[7],mul_out[200][3]);
mul_8x8bit m602 (image[128],filter[8],mul_out[200][4]);

adder_8bit ad66 (mul_out[198][2],mul_out[198][3],mul_out[198][4],mul_out[199][2],mul_out[199][3],mul_out[199][4],mul_out[200][2],mul_out[200][3],mul_out[200][4],conv_out[66]);



mul_8x8bit m603 (image[71],filter[0],mul_out[201][2]);
mul_8x8bit m604 (image[72],filter[1],mul_out[201][3]);
mul_8x8bit m605 (image[73],filter[2],mul_out[201][4]);
mul_8x8bit m606 (image[99],filter[3],mul_out[202][2]);
mul_8x8bit m607 (image[100],filter[4],mul_out[202][3]);
mul_8x8bit m608 (image[101],filter[5],mul_out[202][4]);
mul_8x8bit m609 (image[127],filter[6],mul_out[203][2]);
mul_8x8bit m610 (image[128],filter[7],mul_out[203][3]);
mul_8x8bit m611 (image[129],filter[8],mul_out[203][4]);

adder_8bit ad67 (mul_out[201][2],mul_out[201][3],mul_out[201][4],mul_out[202][2],mul_out[202][3],mul_out[202][4],mul_out[203][2],mul_out[203][3],mul_out[203][4],conv_out[67]);



mul_8x8bit m612 (image[72],filter[0],mul_out[204][2]);
mul_8x8bit m613 (image[73],filter[1],mul_out[204][3]);
mul_8x8bit m614 (image[74],filter[2],mul_out[204][4]);
mul_8x8bit m615 (image[100],filter[3],mul_out[205][2]);
mul_8x8bit m616 (image[101],filter[4],mul_out[205][3]);
mul_8x8bit m617 (image[102],filter[5],mul_out[205][4]);
mul_8x8bit m618 (image[128],filter[6],mul_out[206][2]);
mul_8x8bit m619 (image[129],filter[7],mul_out[206][3]);
mul_8x8bit m620 (image[130],filter[8],mul_out[206][4]);

adder_8bit ad68 (mul_out[204][2],mul_out[204][3],mul_out[204][4],mul_out[205][2],mul_out[205][3],mul_out[205][4],mul_out[206][2],mul_out[206][3],mul_out[206][4],conv_out[68]);



mul_8x8bit m621 (image[73],filter[0],mul_out[207][2]);
mul_8x8bit m622 (image[74],filter[1],mul_out[207][3]);
mul_8x8bit m623 (image[75],filter[2],mul_out[207][4]);
mul_8x8bit m624 (image[101],filter[3],mul_out[208][2]);
mul_8x8bit m625 (image[102],filter[4],mul_out[208][3]);
mul_8x8bit m626 (image[103],filter[5],mul_out[208][4]);
mul_8x8bit m627 (image[129],filter[6],mul_out[209][2]);
mul_8x8bit m628 (image[130],filter[7],mul_out[209][3]);
mul_8x8bit m629 (image[131],filter[8],mul_out[209][4]);

adder_8bit ad69 (mul_out[207][2],mul_out[207][3],mul_out[207][4],mul_out[208][2],mul_out[208][3],mul_out[208][4],mul_out[209][2],mul_out[209][3],mul_out[209][4],conv_out[69]);



mul_8x8bit m630 (image[74],filter[0],mul_out[210][2]);
mul_8x8bit m631 (image[75],filter[1],mul_out[210][3]);
mul_8x8bit m632 (image[76],filter[2],mul_out[210][4]);
mul_8x8bit m633 (image[102],filter[3],mul_out[211][2]);
mul_8x8bit m634 (image[103],filter[4],mul_out[211][3]);
mul_8x8bit m635 (image[104],filter[5],mul_out[211][4]);
mul_8x8bit m636 (image[130],filter[6],mul_out[212][2]);
mul_8x8bit m637 (image[131],filter[7],mul_out[212][3]);
mul_8x8bit m638 (image[132],filter[8],mul_out[212][4]);

adder_8bit ad70 (mul_out[210][2],mul_out[210][3],mul_out[210][4],mul_out[211][2],mul_out[211][3],mul_out[211][4],mul_out[212][2],mul_out[212][3],mul_out[212][4],conv_out[70]);



mul_8x8bit m639 (image[75],filter[0],mul_out[213][2]);
mul_8x8bit m640 (image[76],filter[1],mul_out[213][3]);
mul_8x8bit m641 (image[77],filter[2],mul_out[213][4]);
mul_8x8bit m642 (image[103],filter[3],mul_out[214][2]);
mul_8x8bit m643 (image[104],filter[4],mul_out[214][3]);
mul_8x8bit m644 (image[105],filter[5],mul_out[214][4]);
mul_8x8bit m645 (image[131],filter[6],mul_out[215][2]);
mul_8x8bit m646 (image[132],filter[7],mul_out[215][3]);
mul_8x8bit m647 (image[133],filter[8],mul_out[215][4]);

adder_8bit ad71 (mul_out[213][2],mul_out[213][3],mul_out[213][4],mul_out[214][2],mul_out[214][3],mul_out[214][4],mul_out[215][2],mul_out[215][3],mul_out[215][4],conv_out[71]);



mul_8x8bit m648 (image[76],filter[0],mul_out[216][2]);
mul_8x8bit m649 (image[77],filter[1],mul_out[216][3]);
mul_8x8bit m650 (image[78],filter[2],mul_out[216][4]);
mul_8x8bit m651 (image[104],filter[3],mul_out[217][2]);
mul_8x8bit m652 (image[105],filter[4],mul_out[217][3]);
mul_8x8bit m653 (image[106],filter[5],mul_out[217][4]);
mul_8x8bit m654 (image[132],filter[6],mul_out[218][2]);
mul_8x8bit m655 (image[133],filter[7],mul_out[218][3]);
mul_8x8bit m656 (image[134],filter[8],mul_out[218][4]);

adder_8bit ad72 (mul_out[216][2],mul_out[216][3],mul_out[216][4],mul_out[217][2],mul_out[217][3],mul_out[217][4],mul_out[218][2],mul_out[218][3],mul_out[218][4],conv_out[72]);



mul_8x8bit m657 (image[77],filter[0],mul_out[219][2]);
mul_8x8bit m658 (image[78],filter[1],mul_out[219][3]);
mul_8x8bit m659 (image[79],filter[2],mul_out[219][4]);
mul_8x8bit m660 (image[105],filter[3],mul_out[220][2]);
mul_8x8bit m661 (image[106],filter[4],mul_out[220][3]);
mul_8x8bit m662 (image[107],filter[5],mul_out[220][4]);
mul_8x8bit m663 (image[133],filter[6],mul_out[221][2]);
mul_8x8bit m664 (image[134],filter[7],mul_out[221][3]);
mul_8x8bit m665 (image[135],filter[8],mul_out[221][4]);

adder_8bit ad73 (mul_out[219][2],mul_out[219][3],mul_out[219][4],mul_out[220][2],mul_out[220][3],mul_out[220][4],mul_out[221][2],mul_out[221][3],mul_out[221][4],conv_out[73]);



mul_8x8bit m666 (image[78],filter[0],mul_out[222][2]);
mul_8x8bit m667 (image[79],filter[1],mul_out[222][3]);
mul_8x8bit m668 (image[80],filter[2],mul_out[222][4]);
mul_8x8bit m669 (image[106],filter[3],mul_out[223][2]);
mul_8x8bit m670 (image[107],filter[4],mul_out[223][3]);
mul_8x8bit m671 (image[108],filter[5],mul_out[223][4]);
mul_8x8bit m672 (image[134],filter[6],mul_out[224][2]);
mul_8x8bit m673 (image[135],filter[7],mul_out[224][3]);
mul_8x8bit m674 (image[136],filter[8],mul_out[224][4]);

adder_8bit ad74 (mul_out[222][2],mul_out[222][3],mul_out[222][4],mul_out[223][2],mul_out[223][3],mul_out[223][4],mul_out[224][2],mul_out[224][3],mul_out[224][4],conv_out[74]);



mul_8x8bit m675 (image[79],filter[0],mul_out[225][2]);
mul_8x8bit m676 (image[80],filter[1],mul_out[225][3]);
mul_8x8bit m677 (image[81],filter[2],mul_out[225][4]);
mul_8x8bit m678 (image[107],filter[3],mul_out[226][2]);
mul_8x8bit m679 (image[108],filter[4],mul_out[226][3]);
mul_8x8bit m680 (image[109],filter[5],mul_out[226][4]);
mul_8x8bit m681 (image[135],filter[6],mul_out[227][2]);
mul_8x8bit m682 (image[136],filter[7],mul_out[227][3]);
mul_8x8bit m683 (image[137],filter[8],mul_out[227][4]);

adder_8bit ad75 (mul_out[225][2],mul_out[225][3],mul_out[225][4],mul_out[226][2],mul_out[226][3],mul_out[226][4],mul_out[227][2],mul_out[227][3],mul_out[227][4],conv_out[75]);



mul_8x8bit m684 (image[80],filter[0],mul_out[228][2]);
mul_8x8bit m685 (image[81],filter[1],mul_out[228][3]);
mul_8x8bit m686 (image[82],filter[2],mul_out[228][4]);
mul_8x8bit m687 (image[108],filter[3],mul_out[229][2]);
mul_8x8bit m688 (image[109],filter[4],mul_out[229][3]);
mul_8x8bit m689 (image[110],filter[5],mul_out[229][4]);
mul_8x8bit m690 (image[136],filter[6],mul_out[230][2]);
mul_8x8bit m691 (image[137],filter[7],mul_out[230][3]);
mul_8x8bit m692 (image[138],filter[8],mul_out[230][4]);

adder_8bit ad76 (mul_out[228][2],mul_out[228][3],mul_out[228][4],mul_out[229][2],mul_out[229][3],mul_out[229][4],mul_out[230][2],mul_out[230][3],mul_out[230][4],conv_out[76]);



mul_8x8bit m693 (image[81],filter[0],mul_out[231][2]);
mul_8x8bit m694 (image[82],filter[1],mul_out[231][3]);
mul_8x8bit m695 (image[83],filter[2],mul_out[231][4]);
mul_8x8bit m696 (image[109],filter[3],mul_out[232][2]);
mul_8x8bit m697 (image[110],filter[4],mul_out[232][3]);
mul_8x8bit m698 (image[111],filter[5],mul_out[232][4]);
mul_8x8bit m699 (image[137],filter[6],mul_out[233][2]);
mul_8x8bit m700 (image[138],filter[7],mul_out[233][3]);
mul_8x8bit m701 (image[139],filter[8],mul_out[233][4]);

adder_8bit ad77 (mul_out[231][2],mul_out[231][3],mul_out[231][4],mul_out[232][2],mul_out[232][3],mul_out[232][4],mul_out[233][2],mul_out[233][3],mul_out[233][4],conv_out[77]);



mul_8x8bit m702 (image[84],filter[0],mul_out[234][3]);
mul_8x8bit m703 (image[85],filter[1],mul_out[234][4]);
mul_8x8bit m704 (image[86],filter[2],mul_out[234][5]);
mul_8x8bit m705 (image[112],filter[3],mul_out[235][3]);
mul_8x8bit m706 (image[113],filter[4],mul_out[235][4]);
mul_8x8bit m707 (image[114],filter[5],mul_out[235][5]);
mul_8x8bit m708 (image[140],filter[6],mul_out[236][3]);
mul_8x8bit m709 (image[141],filter[7],mul_out[236][4]);
mul_8x8bit m710 (image[142],filter[8],mul_out[236][5]);

adder_8bit ad78 (mul_out[234][3],mul_out[234][4],mul_out[234][5],mul_out[235][3],mul_out[235][4],mul_out[235][5],mul_out[236][3],mul_out[236][4],mul_out[236][5],conv_out[78]);



mul_8x8bit m711 (image[85],filter[0],mul_out[237][3]);
mul_8x8bit m712 (image[86],filter[1],mul_out[237][4]);
mul_8x8bit m713 (image[87],filter[2],mul_out[237][5]);
mul_8x8bit m714 (image[113],filter[3],mul_out[238][3]);
mul_8x8bit m715 (image[114],filter[4],mul_out[238][4]);
mul_8x8bit m716 (image[115],filter[5],mul_out[238][5]);
mul_8x8bit m717 (image[141],filter[6],mul_out[239][3]);
mul_8x8bit m718 (image[142],filter[7],mul_out[239][4]);
mul_8x8bit m719 (image[143],filter[8],mul_out[239][5]);

adder_8bit ad79 (mul_out[237][3],mul_out[237][4],mul_out[237][5],mul_out[238][3],mul_out[238][4],mul_out[238][5],mul_out[239][3],mul_out[239][4],mul_out[239][5],conv_out[79]);



mul_8x8bit m720 (image[86],filter[0],mul_out[240][3]);
mul_8x8bit m721 (image[87],filter[1],mul_out[240][4]);
mul_8x8bit m722 (image[88],filter[2],mul_out[240][5]);
mul_8x8bit m723 (image[114],filter[3],mul_out[241][3]);
mul_8x8bit m724 (image[115],filter[4],mul_out[241][4]);
mul_8x8bit m725 (image[116],filter[5],mul_out[241][5]);
mul_8x8bit m726 (image[142],filter[6],mul_out[242][3]);
mul_8x8bit m727 (image[143],filter[7],mul_out[242][4]);
mul_8x8bit m728 (image[144],filter[8],mul_out[242][5]);

adder_8bit ad80 (mul_out[240][3],mul_out[240][4],mul_out[240][5],mul_out[241][3],mul_out[241][4],mul_out[241][5],mul_out[242][3],mul_out[242][4],mul_out[242][5],conv_out[80]);



mul_8x8bit m729 (image[87],filter[0],mul_out[243][3]);
mul_8x8bit m730 (image[88],filter[1],mul_out[243][4]);
mul_8x8bit m731 (image[89],filter[2],mul_out[243][5]);
mul_8x8bit m732 (image[115],filter[3],mul_out[244][3]);
mul_8x8bit m733 (image[116],filter[4],mul_out[244][4]);
mul_8x8bit m734 (image[117],filter[5],mul_out[244][5]);
mul_8x8bit m735 (image[143],filter[6],mul_out[245][3]);
mul_8x8bit m736 (image[144],filter[7],mul_out[245][4]);
mul_8x8bit m737 (image[145],filter[8],mul_out[245][5]);

adder_8bit ad81 (mul_out[243][3],mul_out[243][4],mul_out[243][5],mul_out[244][3],mul_out[244][4],mul_out[244][5],mul_out[245][3],mul_out[245][4],mul_out[245][5],conv_out[81]);



mul_8x8bit m738 (image[88],filter[0],mul_out[246][3]);
mul_8x8bit m739 (image[89],filter[1],mul_out[246][4]);
mul_8x8bit m740 (image[90],filter[2],mul_out[246][5]);
mul_8x8bit m741 (image[116],filter[3],mul_out[247][3]);
mul_8x8bit m742 (image[117],filter[4],mul_out[247][4]);
mul_8x8bit m743 (image[118],filter[5],mul_out[247][5]);
mul_8x8bit m744 (image[144],filter[6],mul_out[248][3]);
mul_8x8bit m745 (image[145],filter[7],mul_out[248][4]);
mul_8x8bit m746 (image[146],filter[8],mul_out[248][5]);

adder_8bit ad82 (mul_out[246][3],mul_out[246][4],mul_out[246][5],mul_out[247][3],mul_out[247][4],mul_out[247][5],mul_out[248][3],mul_out[248][4],mul_out[248][5],conv_out[82]);



mul_8x8bit m747 (image[89],filter[0],mul_out[249][3]);
mul_8x8bit m748 (image[90],filter[1],mul_out[249][4]);
mul_8x8bit m749 (image[91],filter[2],mul_out[249][5]);
mul_8x8bit m750 (image[117],filter[3],mul_out[250][3]);
mul_8x8bit m751 (image[118],filter[4],mul_out[250][4]);
mul_8x8bit m752 (image[119],filter[5],mul_out[250][5]);
mul_8x8bit m753 (image[145],filter[6],mul_out[251][3]);
mul_8x8bit m754 (image[146],filter[7],mul_out[251][4]);
mul_8x8bit m755 (image[147],filter[8],mul_out[251][5]);

adder_8bit ad83 (mul_out[249][3],mul_out[249][4],mul_out[249][5],mul_out[250][3],mul_out[250][4],mul_out[250][5],mul_out[251][3],mul_out[251][4],mul_out[251][5],conv_out[83]);



mul_8x8bit m756 (image[90],filter[0],mul_out[252][3]);
mul_8x8bit m757 (image[91],filter[1],mul_out[252][4]);
mul_8x8bit m758 (image[92],filter[2],mul_out[252][5]);
mul_8x8bit m759 (image[118],filter[3],mul_out[253][3]);
mul_8x8bit m760 (image[119],filter[4],mul_out[253][4]);
mul_8x8bit m761 (image[120],filter[5],mul_out[253][5]);
mul_8x8bit m762 (image[146],filter[6],mul_out[254][3]);
mul_8x8bit m763 (image[147],filter[7],mul_out[254][4]);
mul_8x8bit m764 (image[148],filter[8],mul_out[254][5]);

adder_8bit ad84 (mul_out[252][3],mul_out[252][4],mul_out[252][5],mul_out[253][3],mul_out[253][4],mul_out[253][5],mul_out[254][3],mul_out[254][4],mul_out[254][5],conv_out[84]);



mul_8x8bit m765 (image[91],filter[0],mul_out[255][3]);
mul_8x8bit m766 (image[92],filter[1],mul_out[255][4]);
mul_8x8bit m767 (image[93],filter[2],mul_out[255][5]);
mul_8x8bit m768 (image[119],filter[3],mul_out[256][3]);
mul_8x8bit m769 (image[120],filter[4],mul_out[256][4]);
mul_8x8bit m770 (image[121],filter[5],mul_out[256][5]);
mul_8x8bit m771 (image[147],filter[6],mul_out[257][3]);
mul_8x8bit m772 (image[148],filter[7],mul_out[257][4]);
mul_8x8bit m773 (image[149],filter[8],mul_out[257][5]);

adder_8bit ad85 (mul_out[255][3],mul_out[255][4],mul_out[255][5],mul_out[256][3],mul_out[256][4],mul_out[256][5],mul_out[257][3],mul_out[257][4],mul_out[257][5],conv_out[85]);



mul_8x8bit m774 (image[92],filter[0],mul_out[258][3]);
mul_8x8bit m775 (image[93],filter[1],mul_out[258][4]);
mul_8x8bit m776 (image[94],filter[2],mul_out[258][5]);
mul_8x8bit m777 (image[120],filter[3],mul_out[259][3]);
mul_8x8bit m778 (image[121],filter[4],mul_out[259][4]);
mul_8x8bit m779 (image[122],filter[5],mul_out[259][5]);
mul_8x8bit m780 (image[148],filter[6],mul_out[260][3]);
mul_8x8bit m781 (image[149],filter[7],mul_out[260][4]);
mul_8x8bit m782 (image[150],filter[8],mul_out[260][5]);

adder_8bit ad86 (mul_out[258][3],mul_out[258][4],mul_out[258][5],mul_out[259][3],mul_out[259][4],mul_out[259][5],mul_out[260][3],mul_out[260][4],mul_out[260][5],conv_out[86]);



mul_8x8bit m783 (image[93],filter[0],mul_out[261][3]);
mul_8x8bit m784 (image[94],filter[1],mul_out[261][4]);
mul_8x8bit m785 (image[95],filter[2],mul_out[261][5]);
mul_8x8bit m786 (image[121],filter[3],mul_out[262][3]);
mul_8x8bit m787 (image[122],filter[4],mul_out[262][4]);
mul_8x8bit m788 (image[123],filter[5],mul_out[262][5]);
mul_8x8bit m789 (image[149],filter[6],mul_out[263][3]);
mul_8x8bit m790 (image[150],filter[7],mul_out[263][4]);
mul_8x8bit m791 (image[151],filter[8],mul_out[263][5]);

adder_8bit ad87 (mul_out[261][3],mul_out[261][4],mul_out[261][5],mul_out[262][3],mul_out[262][4],mul_out[262][5],mul_out[263][3],mul_out[263][4],mul_out[263][5],conv_out[87]);



mul_8x8bit m792 (image[94],filter[0],mul_out[264][3]);
mul_8x8bit m793 (image[95],filter[1],mul_out[264][4]);
mul_8x8bit m794 (image[96],filter[2],mul_out[264][5]);
mul_8x8bit m795 (image[122],filter[3],mul_out[265][3]);
mul_8x8bit m796 (image[123],filter[4],mul_out[265][4]);
mul_8x8bit m797 (image[124],filter[5],mul_out[265][5]);
mul_8x8bit m798 (image[150],filter[6],mul_out[266][3]);
mul_8x8bit m799 (image[151],filter[7],mul_out[266][4]);
mul_8x8bit m800 (image[152],filter[8],mul_out[266][5]);

adder_8bit ad88 (mul_out[264][3],mul_out[264][4],mul_out[264][5],mul_out[265][3],mul_out[265][4],mul_out[265][5],mul_out[266][3],mul_out[266][4],mul_out[266][5],conv_out[88]);



mul_8x8bit m801 (image[95],filter[0],mul_out[267][3]);
mul_8x8bit m802 (image[96],filter[1],mul_out[267][4]);
mul_8x8bit m803 (image[97],filter[2],mul_out[267][5]);
mul_8x8bit m804 (image[123],filter[3],mul_out[268][3]);
mul_8x8bit m805 (image[124],filter[4],mul_out[268][4]);
mul_8x8bit m806 (image[125],filter[5],mul_out[268][5]);
mul_8x8bit m807 (image[151],filter[6],mul_out[269][3]);
mul_8x8bit m808 (image[152],filter[7],mul_out[269][4]);
mul_8x8bit m809 (image[153],filter[8],mul_out[269][5]);

adder_8bit ad89 (mul_out[267][3],mul_out[267][4],mul_out[267][5],mul_out[268][3],mul_out[268][4],mul_out[268][5],mul_out[269][3],mul_out[269][4],mul_out[269][5],conv_out[89]);



mul_8x8bit m810 (image[96],filter[0],mul_out[270][3]);
mul_8x8bit m811 (image[97],filter[1],mul_out[270][4]);
mul_8x8bit m812 (image[98],filter[2],mul_out[270][5]);
mul_8x8bit m813 (image[124],filter[3],mul_out[271][3]);
mul_8x8bit m814 (image[125],filter[4],mul_out[271][4]);
mul_8x8bit m815 (image[126],filter[5],mul_out[271][5]);
mul_8x8bit m816 (image[152],filter[6],mul_out[272][3]);
mul_8x8bit m817 (image[153],filter[7],mul_out[272][4]);
mul_8x8bit m818 (image[154],filter[8],mul_out[272][5]);

adder_8bit ad90 (mul_out[270][3],mul_out[270][4],mul_out[270][5],mul_out[271][3],mul_out[271][4],mul_out[271][5],mul_out[272][3],mul_out[272][4],mul_out[272][5],conv_out[90]);



mul_8x8bit m819 (image[97],filter[0],mul_out[273][3]);
mul_8x8bit m820 (image[98],filter[1],mul_out[273][4]);
mul_8x8bit m821 (image[99],filter[2],mul_out[273][5]);
mul_8x8bit m822 (image[125],filter[3],mul_out[274][3]);
mul_8x8bit m823 (image[126],filter[4],mul_out[274][4]);
mul_8x8bit m824 (image[127],filter[5],mul_out[274][5]);
mul_8x8bit m825 (image[153],filter[6],mul_out[275][3]);
mul_8x8bit m826 (image[154],filter[7],mul_out[275][4]);
mul_8x8bit m827 (image[155],filter[8],mul_out[275][5]);

adder_8bit ad91 (mul_out[273][3],mul_out[273][4],mul_out[273][5],mul_out[274][3],mul_out[274][4],mul_out[274][5],mul_out[275][3],mul_out[275][4],mul_out[275][5],conv_out[91]);



mul_8x8bit m828 (image[98],filter[0],mul_out[276][3]);
mul_8x8bit m829 (image[99],filter[1],mul_out[276][4]);
mul_8x8bit m830 (image[100],filter[2],mul_out[276][5]);
mul_8x8bit m831 (image[126],filter[3],mul_out[277][3]);
mul_8x8bit m832 (image[127],filter[4],mul_out[277][4]);
mul_8x8bit m833 (image[128],filter[5],mul_out[277][5]);
mul_8x8bit m834 (image[154],filter[6],mul_out[278][3]);
mul_8x8bit m835 (image[155],filter[7],mul_out[278][4]);
mul_8x8bit m836 (image[156],filter[8],mul_out[278][5]);

adder_8bit ad92 (mul_out[276][3],mul_out[276][4],mul_out[276][5],mul_out[277][3],mul_out[277][4],mul_out[277][5],mul_out[278][3],mul_out[278][4],mul_out[278][5],conv_out[92]);



mul_8x8bit m837 (image[99],filter[0],mul_out[279][3]);
mul_8x8bit m838 (image[100],filter[1],mul_out[279][4]);
mul_8x8bit m839 (image[101],filter[2],mul_out[279][5]);
mul_8x8bit m840 (image[127],filter[3],mul_out[280][3]);
mul_8x8bit m841 (image[128],filter[4],mul_out[280][4]);
mul_8x8bit m842 (image[129],filter[5],mul_out[280][5]);
mul_8x8bit m843 (image[155],filter[6],mul_out[281][3]);
mul_8x8bit m844 (image[156],filter[7],mul_out[281][4]);
mul_8x8bit m845 (image[157],filter[8],mul_out[281][5]);

adder_8bit ad93 (mul_out[279][3],mul_out[279][4],mul_out[279][5],mul_out[280][3],mul_out[280][4],mul_out[280][5],mul_out[281][3],mul_out[281][4],mul_out[281][5],conv_out[93]);



mul_8x8bit m846 (image[100],filter[0],mul_out[282][3]);
mul_8x8bit m847 (image[101],filter[1],mul_out[282][4]);
mul_8x8bit m848 (image[102],filter[2],mul_out[282][5]);
mul_8x8bit m849 (image[128],filter[3],mul_out[283][3]);
mul_8x8bit m850 (image[129],filter[4],mul_out[283][4]);
mul_8x8bit m851 (image[130],filter[5],mul_out[283][5]);
mul_8x8bit m852 (image[156],filter[6],mul_out[284][3]);
mul_8x8bit m853 (image[157],filter[7],mul_out[284][4]);
mul_8x8bit m854 (image[158],filter[8],mul_out[284][5]);

adder_8bit ad94 (mul_out[282][3],mul_out[282][4],mul_out[282][5],mul_out[283][3],mul_out[283][4],mul_out[283][5],mul_out[284][3],mul_out[284][4],mul_out[284][5],conv_out[94]);



mul_8x8bit m855 (image[101],filter[0],mul_out[285][3]);
mul_8x8bit m856 (image[102],filter[1],mul_out[285][4]);
mul_8x8bit m857 (image[103],filter[2],mul_out[285][5]);
mul_8x8bit m858 (image[129],filter[3],mul_out[286][3]);
mul_8x8bit m859 (image[130],filter[4],mul_out[286][4]);
mul_8x8bit m860 (image[131],filter[5],mul_out[286][5]);
mul_8x8bit m861 (image[157],filter[6],mul_out[287][3]);
mul_8x8bit m862 (image[158],filter[7],mul_out[287][4]);
mul_8x8bit m863 (image[159],filter[8],mul_out[287][5]);

adder_8bit ad95 (mul_out[285][3],mul_out[285][4],mul_out[285][5],mul_out[286][3],mul_out[286][4],mul_out[286][5],mul_out[287][3],mul_out[287][4],mul_out[287][5],conv_out[95]);



mul_8x8bit m864 (image[102],filter[0],mul_out[288][3]);
mul_8x8bit m865 (image[103],filter[1],mul_out[288][4]);
mul_8x8bit m866 (image[104],filter[2],mul_out[288][5]);
mul_8x8bit m867 (image[130],filter[3],mul_out[289][3]);
mul_8x8bit m868 (image[131],filter[4],mul_out[289][4]);
mul_8x8bit m869 (image[132],filter[5],mul_out[289][5]);
mul_8x8bit m870 (image[158],filter[6],mul_out[290][3]);
mul_8x8bit m871 (image[159],filter[7],mul_out[290][4]);
mul_8x8bit m872 (image[160],filter[8],mul_out[290][5]);

adder_8bit ad96 (mul_out[288][3],mul_out[288][4],mul_out[288][5],mul_out[289][3],mul_out[289][4],mul_out[289][5],mul_out[290][3],mul_out[290][4],mul_out[290][5],conv_out[96]);



mul_8x8bit m873 (image[103],filter[0],mul_out[291][3]);
mul_8x8bit m874 (image[104],filter[1],mul_out[291][4]);
mul_8x8bit m875 (image[105],filter[2],mul_out[291][5]);
mul_8x8bit m876 (image[131],filter[3],mul_out[292][3]);
mul_8x8bit m877 (image[132],filter[4],mul_out[292][4]);
mul_8x8bit m878 (image[133],filter[5],mul_out[292][5]);
mul_8x8bit m879 (image[159],filter[6],mul_out[293][3]);
mul_8x8bit m880 (image[160],filter[7],mul_out[293][4]);
mul_8x8bit m881 (image[161],filter[8],mul_out[293][5]);

adder_8bit ad97 (mul_out[291][3],mul_out[291][4],mul_out[291][5],mul_out[292][3],mul_out[292][4],mul_out[292][5],mul_out[293][3],mul_out[293][4],mul_out[293][5],conv_out[97]);



mul_8x8bit m882 (image[104],filter[0],mul_out[294][3]);
mul_8x8bit m883 (image[105],filter[1],mul_out[294][4]);
mul_8x8bit m884 (image[106],filter[2],mul_out[294][5]);
mul_8x8bit m885 (image[132],filter[3],mul_out[295][3]);
mul_8x8bit m886 (image[133],filter[4],mul_out[295][4]);
mul_8x8bit m887 (image[134],filter[5],mul_out[295][5]);
mul_8x8bit m888 (image[160],filter[6],mul_out[296][3]);
mul_8x8bit m889 (image[161],filter[7],mul_out[296][4]);
mul_8x8bit m890 (image[162],filter[8],mul_out[296][5]);

adder_8bit ad98 (mul_out[294][3],mul_out[294][4],mul_out[294][5],mul_out[295][3],mul_out[295][4],mul_out[295][5],mul_out[296][3],mul_out[296][4],mul_out[296][5],conv_out[98]);



mul_8x8bit m891 (image[105],filter[0],mul_out[297][3]);
mul_8x8bit m892 (image[106],filter[1],mul_out[297][4]);
mul_8x8bit m893 (image[107],filter[2],mul_out[297][5]);
mul_8x8bit m894 (image[133],filter[3],mul_out[298][3]);
mul_8x8bit m895 (image[134],filter[4],mul_out[298][4]);
mul_8x8bit m896 (image[135],filter[5],mul_out[298][5]);
mul_8x8bit m897 (image[161],filter[6],mul_out[299][3]);
mul_8x8bit m898 (image[162],filter[7],mul_out[299][4]);
mul_8x8bit m899 (image[163],filter[8],mul_out[299][5]);

adder_8bit ad99 (mul_out[297][3],mul_out[297][4],mul_out[297][5],mul_out[298][3],mul_out[298][4],mul_out[298][5],mul_out[299][3],mul_out[299][4],mul_out[299][5],conv_out[99]);



mul_8x8bit m900 (image[106],filter[0],mul_out[300][3]);
mul_8x8bit m901 (image[107],filter[1],mul_out[300][4]);
mul_8x8bit m902 (image[108],filter[2],mul_out[300][5]);
mul_8x8bit m903 (image[134],filter[3],mul_out[301][3]);
mul_8x8bit m904 (image[135],filter[4],mul_out[301][4]);
mul_8x8bit m905 (image[136],filter[5],mul_out[301][5]);
mul_8x8bit m906 (image[162],filter[6],mul_out[302][3]);
mul_8x8bit m907 (image[163],filter[7],mul_out[302][4]);
mul_8x8bit m908 (image[164],filter[8],mul_out[302][5]);

adder_8bit ad100 (mul_out[300][3],mul_out[300][4],mul_out[300][5],mul_out[301][3],mul_out[301][4],mul_out[301][5],mul_out[302][3],mul_out[302][4],mul_out[302][5],conv_out[100]);



mul_8x8bit m909 (image[107],filter[0],mul_out[303][3]);
mul_8x8bit m910 (image[108],filter[1],mul_out[303][4]);
mul_8x8bit m911 (image[109],filter[2],mul_out[303][5]);
mul_8x8bit m912 (image[135],filter[3],mul_out[304][3]);
mul_8x8bit m913 (image[136],filter[4],mul_out[304][4]);
mul_8x8bit m914 (image[137],filter[5],mul_out[304][5]);
mul_8x8bit m915 (image[163],filter[6],mul_out[305][3]);
mul_8x8bit m916 (image[164],filter[7],mul_out[305][4]);
mul_8x8bit m917 (image[165],filter[8],mul_out[305][5]);

adder_8bit ad101 (mul_out[303][3],mul_out[303][4],mul_out[303][5],mul_out[304][3],mul_out[304][4],mul_out[304][5],mul_out[305][3],mul_out[305][4],mul_out[305][5],conv_out[101]);



mul_8x8bit m918 (image[108],filter[0],mul_out[306][3]);
mul_8x8bit m919 (image[109],filter[1],mul_out[306][4]);
mul_8x8bit m920 (image[110],filter[2],mul_out[306][5]);
mul_8x8bit m921 (image[136],filter[3],mul_out[307][3]);
mul_8x8bit m922 (image[137],filter[4],mul_out[307][4]);
mul_8x8bit m923 (image[138],filter[5],mul_out[307][5]);
mul_8x8bit m924 (image[164],filter[6],mul_out[308][3]);
mul_8x8bit m925 (image[165],filter[7],mul_out[308][4]);
mul_8x8bit m926 (image[166],filter[8],mul_out[308][5]);

adder_8bit ad102 (mul_out[306][3],mul_out[306][4],mul_out[306][5],mul_out[307][3],mul_out[307][4],mul_out[307][5],mul_out[308][3],mul_out[308][4],mul_out[308][5],conv_out[102]);



mul_8x8bit m927 (image[109],filter[0],mul_out[309][3]);
mul_8x8bit m928 (image[110],filter[1],mul_out[309][4]);
mul_8x8bit m929 (image[111],filter[2],mul_out[309][5]);
mul_8x8bit m930 (image[137],filter[3],mul_out[310][3]);
mul_8x8bit m931 (image[138],filter[4],mul_out[310][4]);
mul_8x8bit m932 (image[139],filter[5],mul_out[310][5]);
mul_8x8bit m933 (image[165],filter[6],mul_out[311][3]);
mul_8x8bit m934 (image[166],filter[7],mul_out[311][4]);
mul_8x8bit m935 (image[167],filter[8],mul_out[311][5]);

adder_8bit ad103 (mul_out[309][3],mul_out[309][4],mul_out[309][5],mul_out[310][3],mul_out[310][4],mul_out[310][5],mul_out[311][3],mul_out[311][4],mul_out[311][5],conv_out[103]);



mul_8x8bit m936 (image[112],filter[0],mul_out[312][4]);
mul_8x8bit m937 (image[113],filter[1],mul_out[312][5]);
mul_8x8bit m938 (image[114],filter[2],mul_out[312][6]);
mul_8x8bit m939 (image[140],filter[3],mul_out[313][4]);
mul_8x8bit m940 (image[141],filter[4],mul_out[313][5]);
mul_8x8bit m941 (image[142],filter[5],mul_out[313][6]);
mul_8x8bit m942 (image[168],filter[6],mul_out[314][4]);
mul_8x8bit m943 (image[169],filter[7],mul_out[314][5]);
mul_8x8bit m944 (image[170],filter[8],mul_out[314][6]);

adder_8bit ad104 (mul_out[312][4],mul_out[312][5],mul_out[312][6],mul_out[313][4],mul_out[313][5],mul_out[313][6],mul_out[314][4],mul_out[314][5],mul_out[314][6],conv_out[104]);



mul_8x8bit m945 (image[113],filter[0],mul_out[315][4]);
mul_8x8bit m946 (image[114],filter[1],mul_out[315][5]);
mul_8x8bit m947 (image[115],filter[2],mul_out[315][6]);
mul_8x8bit m948 (image[141],filter[3],mul_out[316][4]);
mul_8x8bit m949 (image[142],filter[4],mul_out[316][5]);
mul_8x8bit m950 (image[143],filter[5],mul_out[316][6]);
mul_8x8bit m951 (image[169],filter[6],mul_out[317][4]);
mul_8x8bit m952 (image[170],filter[7],mul_out[317][5]);
mul_8x8bit m953 (image[171],filter[8],mul_out[317][6]);

adder_8bit ad105 (mul_out[315][4],mul_out[315][5],mul_out[315][6],mul_out[316][4],mul_out[316][5],mul_out[316][6],mul_out[317][4],mul_out[317][5],mul_out[317][6],conv_out[105]);



mul_8x8bit m954 (image[114],filter[0],mul_out[318][4]);
mul_8x8bit m955 (image[115],filter[1],mul_out[318][5]);
mul_8x8bit m956 (image[116],filter[2],mul_out[318][6]);
mul_8x8bit m957 (image[142],filter[3],mul_out[319][4]);
mul_8x8bit m958 (image[143],filter[4],mul_out[319][5]);
mul_8x8bit m959 (image[144],filter[5],mul_out[319][6]);
mul_8x8bit m960 (image[170],filter[6],mul_out[320][4]);
mul_8x8bit m961 (image[171],filter[7],mul_out[320][5]);
mul_8x8bit m962 (image[172],filter[8],mul_out[320][6]);

adder_8bit ad106 (mul_out[318][4],mul_out[318][5],mul_out[318][6],mul_out[319][4],mul_out[319][5],mul_out[319][6],mul_out[320][4],mul_out[320][5],mul_out[320][6],conv_out[106]);



mul_8x8bit m963 (image[115],filter[0],mul_out[321][4]);
mul_8x8bit m964 (image[116],filter[1],mul_out[321][5]);
mul_8x8bit m965 (image[117],filter[2],mul_out[321][6]);
mul_8x8bit m966 (image[143],filter[3],mul_out[322][4]);
mul_8x8bit m967 (image[144],filter[4],mul_out[322][5]);
mul_8x8bit m968 (image[145],filter[5],mul_out[322][6]);
mul_8x8bit m969 (image[171],filter[6],mul_out[323][4]);
mul_8x8bit m970 (image[172],filter[7],mul_out[323][5]);
mul_8x8bit m971 (image[173],filter[8],mul_out[323][6]);

adder_8bit ad107 (mul_out[321][4],mul_out[321][5],mul_out[321][6],mul_out[322][4],mul_out[322][5],mul_out[322][6],mul_out[323][4],mul_out[323][5],mul_out[323][6],conv_out[107]);



mul_8x8bit m972 (image[116],filter[0],mul_out[324][4]);
mul_8x8bit m973 (image[117],filter[1],mul_out[324][5]);
mul_8x8bit m974 (image[118],filter[2],mul_out[324][6]);
mul_8x8bit m975 (image[144],filter[3],mul_out[325][4]);
mul_8x8bit m976 (image[145],filter[4],mul_out[325][5]);
mul_8x8bit m977 (image[146],filter[5],mul_out[325][6]);
mul_8x8bit m978 (image[172],filter[6],mul_out[326][4]);
mul_8x8bit m979 (image[173],filter[7],mul_out[326][5]);
mul_8x8bit m980 (image[174],filter[8],mul_out[326][6]);

adder_8bit ad108 (mul_out[324][4],mul_out[324][5],mul_out[324][6],mul_out[325][4],mul_out[325][5],mul_out[325][6],mul_out[326][4],mul_out[326][5],mul_out[326][6],conv_out[108]);



mul_8x8bit m981 (image[117],filter[0],mul_out[327][4]);
mul_8x8bit m982 (image[118],filter[1],mul_out[327][5]);
mul_8x8bit m983 (image[119],filter[2],mul_out[327][6]);
mul_8x8bit m984 (image[145],filter[3],mul_out[328][4]);
mul_8x8bit m985 (image[146],filter[4],mul_out[328][5]);
mul_8x8bit m986 (image[147],filter[5],mul_out[328][6]);
mul_8x8bit m987 (image[173],filter[6],mul_out[329][4]);
mul_8x8bit m988 (image[174],filter[7],mul_out[329][5]);
mul_8x8bit m989 (image[175],filter[8],mul_out[329][6]);

adder_8bit ad109 (mul_out[327][4],mul_out[327][5],mul_out[327][6],mul_out[328][4],mul_out[328][5],mul_out[328][6],mul_out[329][4],mul_out[329][5],mul_out[329][6],conv_out[109]);



mul_8x8bit m990 (image[118],filter[0],mul_out[330][4]);
mul_8x8bit m991 (image[119],filter[1],mul_out[330][5]);
mul_8x8bit m992 (image[120],filter[2],mul_out[330][6]);
mul_8x8bit m993 (image[146],filter[3],mul_out[331][4]);
mul_8x8bit m994 (image[147],filter[4],mul_out[331][5]);
mul_8x8bit m995 (image[148],filter[5],mul_out[331][6]);
mul_8x8bit m996 (image[174],filter[6],mul_out[332][4]);
mul_8x8bit m997 (image[175],filter[7],mul_out[332][5]);
mul_8x8bit m998 (image[176],filter[8],mul_out[332][6]);

adder_8bit ad110 (mul_out[330][4],mul_out[330][5],mul_out[330][6],mul_out[331][4],mul_out[331][5],mul_out[331][6],mul_out[332][4],mul_out[332][5],mul_out[332][6],conv_out[110]);



mul_8x8bit m999 (image[119],filter[0],mul_out[333][4]);
mul_8x8bit m1000 (image[120],filter[1],mul_out[333][5]);
mul_8x8bit m1001 (image[121],filter[2],mul_out[333][6]);
mul_8x8bit m1002 (image[147],filter[3],mul_out[334][4]);
mul_8x8bit m1003 (image[148],filter[4],mul_out[334][5]);
mul_8x8bit m1004 (image[149],filter[5],mul_out[334][6]);
mul_8x8bit m1005 (image[175],filter[6],mul_out[335][4]);
mul_8x8bit m1006 (image[176],filter[7],mul_out[335][5]);
mul_8x8bit m1007 (image[177],filter[8],mul_out[335][6]);

adder_8bit ad111 (mul_out[333][4],mul_out[333][5],mul_out[333][6],mul_out[334][4],mul_out[334][5],mul_out[334][6],mul_out[335][4],mul_out[335][5],mul_out[335][6],conv_out[111]);



mul_8x8bit m1008 (image[120],filter[0],mul_out[336][4]);
mul_8x8bit m1009 (image[121],filter[1],mul_out[336][5]);
mul_8x8bit m1010 (image[122],filter[2],mul_out[336][6]);
mul_8x8bit m1011 (image[148],filter[3],mul_out[337][4]);
mul_8x8bit m1012 (image[149],filter[4],mul_out[337][5]);
mul_8x8bit m1013 (image[150],filter[5],mul_out[337][6]);
mul_8x8bit m1014 (image[176],filter[6],mul_out[338][4]);
mul_8x8bit m1015 (image[177],filter[7],mul_out[338][5]);
mul_8x8bit m1016 (image[178],filter[8],mul_out[338][6]);

adder_8bit ad112 (mul_out[336][4],mul_out[336][5],mul_out[336][6],mul_out[337][4],mul_out[337][5],mul_out[337][6],mul_out[338][4],mul_out[338][5],mul_out[338][6],conv_out[112]);



mul_8x8bit m1017 (image[121],filter[0],mul_out[339][4]);
mul_8x8bit m1018 (image[122],filter[1],mul_out[339][5]);
mul_8x8bit m1019 (image[123],filter[2],mul_out[339][6]);
mul_8x8bit m1020 (image[149],filter[3],mul_out[340][4]);
mul_8x8bit m1021 (image[150],filter[4],mul_out[340][5]);
mul_8x8bit m1022 (image[151],filter[5],mul_out[340][6]);
mul_8x8bit m1023 (image[177],filter[6],mul_out[341][4]);
mul_8x8bit m1024 (image[178],filter[7],mul_out[341][5]);
mul_8x8bit m1025 (image[179],filter[8],mul_out[341][6]);

adder_8bit ad113 (mul_out[339][4],mul_out[339][5],mul_out[339][6],mul_out[340][4],mul_out[340][5],mul_out[340][6],mul_out[341][4],mul_out[341][5],mul_out[341][6],conv_out[113]);



mul_8x8bit m1026 (image[122],filter[0],mul_out[342][4]);
mul_8x8bit m1027 (image[123],filter[1],mul_out[342][5]);
mul_8x8bit m1028 (image[124],filter[2],mul_out[342][6]);
mul_8x8bit m1029 (image[150],filter[3],mul_out[343][4]);
mul_8x8bit m1030 (image[151],filter[4],mul_out[343][5]);
mul_8x8bit m1031 (image[152],filter[5],mul_out[343][6]);
mul_8x8bit m1032 (image[178],filter[6],mul_out[344][4]);
mul_8x8bit m1033 (image[179],filter[7],mul_out[344][5]);
mul_8x8bit m1034 (image[180],filter[8],mul_out[344][6]);

adder_8bit ad114 (mul_out[342][4],mul_out[342][5],mul_out[342][6],mul_out[343][4],mul_out[343][5],mul_out[343][6],mul_out[344][4],mul_out[344][5],mul_out[344][6],conv_out[114]);



mul_8x8bit m1035 (image[123],filter[0],mul_out[345][4]);
mul_8x8bit m1036 (image[124],filter[1],mul_out[345][5]);
mul_8x8bit m1037 (image[125],filter[2],mul_out[345][6]);
mul_8x8bit m1038 (image[151],filter[3],mul_out[346][4]);
mul_8x8bit m1039 (image[152],filter[4],mul_out[346][5]);
mul_8x8bit m1040 (image[153],filter[5],mul_out[346][6]);
mul_8x8bit m1041 (image[179],filter[6],mul_out[347][4]);
mul_8x8bit m1042 (image[180],filter[7],mul_out[347][5]);
mul_8x8bit m1043 (image[181],filter[8],mul_out[347][6]);

adder_8bit ad115 (mul_out[345][4],mul_out[345][5],mul_out[345][6],mul_out[346][4],mul_out[346][5],mul_out[346][6],mul_out[347][4],mul_out[347][5],mul_out[347][6],conv_out[115]);



mul_8x8bit m1044 (image[124],filter[0],mul_out[348][4]);
mul_8x8bit m1045 (image[125],filter[1],mul_out[348][5]);
mul_8x8bit m1046 (image[126],filter[2],mul_out[348][6]);
mul_8x8bit m1047 (image[152],filter[3],mul_out[349][4]);
mul_8x8bit m1048 (image[153],filter[4],mul_out[349][5]);
mul_8x8bit m1049 (image[154],filter[5],mul_out[349][6]);
mul_8x8bit m1050 (image[180],filter[6],mul_out[350][4]);
mul_8x8bit m1051 (image[181],filter[7],mul_out[350][5]);
mul_8x8bit m1052 (image[182],filter[8],mul_out[350][6]);

adder_8bit ad116 (mul_out[348][4],mul_out[348][5],mul_out[348][6],mul_out[349][4],mul_out[349][5],mul_out[349][6],mul_out[350][4],mul_out[350][5],mul_out[350][6],conv_out[116]);



mul_8x8bit m1053 (image[125],filter[0],mul_out[351][4]);
mul_8x8bit m1054 (image[126],filter[1],mul_out[351][5]);
mul_8x8bit m1055 (image[127],filter[2],mul_out[351][6]);
mul_8x8bit m1056 (image[153],filter[3],mul_out[352][4]);
mul_8x8bit m1057 (image[154],filter[4],mul_out[352][5]);
mul_8x8bit m1058 (image[155],filter[5],mul_out[352][6]);
mul_8x8bit m1059 (image[181],filter[6],mul_out[353][4]);
mul_8x8bit m1060 (image[182],filter[7],mul_out[353][5]);
mul_8x8bit m1061 (image[183],filter[8],mul_out[353][6]);

adder_8bit ad117 (mul_out[351][4],mul_out[351][5],mul_out[351][6],mul_out[352][4],mul_out[352][5],mul_out[352][6],mul_out[353][4],mul_out[353][5],mul_out[353][6],conv_out[117]);



mul_8x8bit m1062 (image[126],filter[0],mul_out[354][4]);
mul_8x8bit m1063 (image[127],filter[1],mul_out[354][5]);
mul_8x8bit m1064 (image[128],filter[2],mul_out[354][6]);
mul_8x8bit m1065 (image[154],filter[3],mul_out[355][4]);
mul_8x8bit m1066 (image[155],filter[4],mul_out[355][5]);
mul_8x8bit m1067 (image[156],filter[5],mul_out[355][6]);
mul_8x8bit m1068 (image[182],filter[6],mul_out[356][4]);
mul_8x8bit m1069 (image[183],filter[7],mul_out[356][5]);
mul_8x8bit m1070 (image[184],filter[8],mul_out[356][6]);

adder_8bit ad118 (mul_out[354][4],mul_out[354][5],mul_out[354][6],mul_out[355][4],mul_out[355][5],mul_out[355][6],mul_out[356][4],mul_out[356][5],mul_out[356][6],conv_out[118]);



mul_8x8bit m1071 (image[127],filter[0],mul_out[357][4]);
mul_8x8bit m1072 (image[128],filter[1],mul_out[357][5]);
mul_8x8bit m1073 (image[129],filter[2],mul_out[357][6]);
mul_8x8bit m1074 (image[155],filter[3],mul_out[358][4]);
mul_8x8bit m1075 (image[156],filter[4],mul_out[358][5]);
mul_8x8bit m1076 (image[157],filter[5],mul_out[358][6]);
mul_8x8bit m1077 (image[183],filter[6],mul_out[359][4]);
mul_8x8bit m1078 (image[184],filter[7],mul_out[359][5]);
mul_8x8bit m1079 (image[185],filter[8],mul_out[359][6]);

adder_8bit ad119 (mul_out[357][4],mul_out[357][5],mul_out[357][6],mul_out[358][4],mul_out[358][5],mul_out[358][6],mul_out[359][4],mul_out[359][5],mul_out[359][6],conv_out[119]);



mul_8x8bit m1080 (image[128],filter[0],mul_out[360][4]);
mul_8x8bit m1081 (image[129],filter[1],mul_out[360][5]);
mul_8x8bit m1082 (image[130],filter[2],mul_out[360][6]);
mul_8x8bit m1083 (image[156],filter[3],mul_out[361][4]);
mul_8x8bit m1084 (image[157],filter[4],mul_out[361][5]);
mul_8x8bit m1085 (image[158],filter[5],mul_out[361][6]);
mul_8x8bit m1086 (image[184],filter[6],mul_out[362][4]);
mul_8x8bit m1087 (image[185],filter[7],mul_out[362][5]);
mul_8x8bit m1088 (image[186],filter[8],mul_out[362][6]);

adder_8bit ad120 (mul_out[360][4],mul_out[360][5],mul_out[360][6],mul_out[361][4],mul_out[361][5],mul_out[361][6],mul_out[362][4],mul_out[362][5],mul_out[362][6],conv_out[120]);



mul_8x8bit m1089 (image[129],filter[0],mul_out[363][4]);
mul_8x8bit m1090 (image[130],filter[1],mul_out[363][5]);
mul_8x8bit m1091 (image[131],filter[2],mul_out[363][6]);
mul_8x8bit m1092 (image[157],filter[3],mul_out[364][4]);
mul_8x8bit m1093 (image[158],filter[4],mul_out[364][5]);
mul_8x8bit m1094 (image[159],filter[5],mul_out[364][6]);
mul_8x8bit m1095 (image[185],filter[6],mul_out[365][4]);
mul_8x8bit m1096 (image[186],filter[7],mul_out[365][5]);
mul_8x8bit m1097 (image[187],filter[8],mul_out[365][6]);

adder_8bit ad121 (mul_out[363][4],mul_out[363][5],mul_out[363][6],mul_out[364][4],mul_out[364][5],mul_out[364][6],mul_out[365][4],mul_out[365][5],mul_out[365][6],conv_out[121]);



mul_8x8bit m1098 (image[130],filter[0],mul_out[366][4]);
mul_8x8bit m1099 (image[131],filter[1],mul_out[366][5]);
mul_8x8bit m1100 (image[132],filter[2],mul_out[366][6]);
mul_8x8bit m1101 (image[158],filter[3],mul_out[367][4]);
mul_8x8bit m1102 (image[159],filter[4],mul_out[367][5]);
mul_8x8bit m1103 (image[160],filter[5],mul_out[367][6]);
mul_8x8bit m1104 (image[186],filter[6],mul_out[368][4]);
mul_8x8bit m1105 (image[187],filter[7],mul_out[368][5]);
mul_8x8bit m1106 (image[188],filter[8],mul_out[368][6]);

adder_8bit ad122 (mul_out[366][4],mul_out[366][5],mul_out[366][6],mul_out[367][4],mul_out[367][5],mul_out[367][6],mul_out[368][4],mul_out[368][5],mul_out[368][6],conv_out[122]);



mul_8x8bit m1107 (image[131],filter[0],mul_out[369][4]);
mul_8x8bit m1108 (image[132],filter[1],mul_out[369][5]);
mul_8x8bit m1109 (image[133],filter[2],mul_out[369][6]);
mul_8x8bit m1110 (image[159],filter[3],mul_out[370][4]);
mul_8x8bit m1111 (image[160],filter[4],mul_out[370][5]);
mul_8x8bit m1112 (image[161],filter[5],mul_out[370][6]);
mul_8x8bit m1113 (image[187],filter[6],mul_out[371][4]);
mul_8x8bit m1114 (image[188],filter[7],mul_out[371][5]);
mul_8x8bit m1115 (image[189],filter[8],mul_out[371][6]);

adder_8bit ad123 (mul_out[369][4],mul_out[369][5],mul_out[369][6],mul_out[370][4],mul_out[370][5],mul_out[370][6],mul_out[371][4],mul_out[371][5],mul_out[371][6],conv_out[123]);



mul_8x8bit m1116 (image[132],filter[0],mul_out[372][4]);
mul_8x8bit m1117 (image[133],filter[1],mul_out[372][5]);
mul_8x8bit m1118 (image[134],filter[2],mul_out[372][6]);
mul_8x8bit m1119 (image[160],filter[3],mul_out[373][4]);
mul_8x8bit m1120 (image[161],filter[4],mul_out[373][5]);
mul_8x8bit m1121 (image[162],filter[5],mul_out[373][6]);
mul_8x8bit m1122 (image[188],filter[6],mul_out[374][4]);
mul_8x8bit m1123 (image[189],filter[7],mul_out[374][5]);
mul_8x8bit m1124 (image[190],filter[8],mul_out[374][6]);

adder_8bit ad124 (mul_out[372][4],mul_out[372][5],mul_out[372][6],mul_out[373][4],mul_out[373][5],mul_out[373][6],mul_out[374][4],mul_out[374][5],mul_out[374][6],conv_out[124]);



mul_8x8bit m1125 (image[133],filter[0],mul_out[375][4]);
mul_8x8bit m1126 (image[134],filter[1],mul_out[375][5]);
mul_8x8bit m1127 (image[135],filter[2],mul_out[375][6]);
mul_8x8bit m1128 (image[161],filter[3],mul_out[376][4]);
mul_8x8bit m1129 (image[162],filter[4],mul_out[376][5]);
mul_8x8bit m1130 (image[163],filter[5],mul_out[376][6]);
mul_8x8bit m1131 (image[189],filter[6],mul_out[377][4]);
mul_8x8bit m1132 (image[190],filter[7],mul_out[377][5]);
mul_8x8bit m1133 (image[191],filter[8],mul_out[377][6]);

adder_8bit ad125 (mul_out[375][4],mul_out[375][5],mul_out[375][6],mul_out[376][4],mul_out[376][5],mul_out[376][6],mul_out[377][4],mul_out[377][5],mul_out[377][6],conv_out[125]);



mul_8x8bit m1134 (image[134],filter[0],mul_out[378][4]);
mul_8x8bit m1135 (image[135],filter[1],mul_out[378][5]);
mul_8x8bit m1136 (image[136],filter[2],mul_out[378][6]);
mul_8x8bit m1137 (image[162],filter[3],mul_out[379][4]);
mul_8x8bit m1138 (image[163],filter[4],mul_out[379][5]);
mul_8x8bit m1139 (image[164],filter[5],mul_out[379][6]);
mul_8x8bit m1140 (image[190],filter[6],mul_out[380][4]);
mul_8x8bit m1141 (image[191],filter[7],mul_out[380][5]);
mul_8x8bit m1142 (image[192],filter[8],mul_out[380][6]);

adder_8bit ad126 (mul_out[378][4],mul_out[378][5],mul_out[378][6],mul_out[379][4],mul_out[379][5],mul_out[379][6],mul_out[380][4],mul_out[380][5],mul_out[380][6],conv_out[126]);



mul_8x8bit m1143 (image[135],filter[0],mul_out[381][4]);
mul_8x8bit m1144 (image[136],filter[1],mul_out[381][5]);
mul_8x8bit m1145 (image[137],filter[2],mul_out[381][6]);
mul_8x8bit m1146 (image[163],filter[3],mul_out[382][4]);
mul_8x8bit m1147 (image[164],filter[4],mul_out[382][5]);
mul_8x8bit m1148 (image[165],filter[5],mul_out[382][6]);
mul_8x8bit m1149 (image[191],filter[6],mul_out[383][4]);
mul_8x8bit m1150 (image[192],filter[7],mul_out[383][5]);
mul_8x8bit m1151 (image[193],filter[8],mul_out[383][6]);

adder_8bit ad127 (mul_out[381][4],mul_out[381][5],mul_out[381][6],mul_out[382][4],mul_out[382][5],mul_out[382][6],mul_out[383][4],mul_out[383][5],mul_out[383][6],conv_out[127]);



mul_8x8bit m1152 (image[136],filter[0],mul_out[384][4]);
mul_8x8bit m1153 (image[137],filter[1],mul_out[384][5]);
mul_8x8bit m1154 (image[138],filter[2],mul_out[384][6]);
mul_8x8bit m1155 (image[164],filter[3],mul_out[385][4]);
mul_8x8bit m1156 (image[165],filter[4],mul_out[385][5]);
mul_8x8bit m1157 (image[166],filter[5],mul_out[385][6]);
mul_8x8bit m1158 (image[192],filter[6],mul_out[386][4]);
mul_8x8bit m1159 (image[193],filter[7],mul_out[386][5]);
mul_8x8bit m1160 (image[194],filter[8],mul_out[386][6]);

adder_8bit ad128 (mul_out[384][4],mul_out[384][5],mul_out[384][6],mul_out[385][4],mul_out[385][5],mul_out[385][6],mul_out[386][4],mul_out[386][5],mul_out[386][6],conv_out[128]);



mul_8x8bit m1161 (image[137],filter[0],mul_out[387][4]);
mul_8x8bit m1162 (image[138],filter[1],mul_out[387][5]);
mul_8x8bit m1163 (image[139],filter[2],mul_out[387][6]);
mul_8x8bit m1164 (image[165],filter[3],mul_out[388][4]);
mul_8x8bit m1165 (image[166],filter[4],mul_out[388][5]);
mul_8x8bit m1166 (image[167],filter[5],mul_out[388][6]);
mul_8x8bit m1167 (image[193],filter[6],mul_out[389][4]);
mul_8x8bit m1168 (image[194],filter[7],mul_out[389][5]);
mul_8x8bit m1169 (image[195],filter[8],mul_out[389][6]);

adder_8bit ad129 (mul_out[387][4],mul_out[387][5],mul_out[387][6],mul_out[388][4],mul_out[388][5],mul_out[388][6],mul_out[389][4],mul_out[389][5],mul_out[389][6],conv_out[129]);



mul_8x8bit m1170 (image[140],filter[0],mul_out[390][5]);
mul_8x8bit m1171 (image[141],filter[1],mul_out[390][6]);
mul_8x8bit m1172 (image[142],filter[2],mul_out[390][7]);
mul_8x8bit m1173 (image[168],filter[3],mul_out[391][5]);
mul_8x8bit m1174 (image[169],filter[4],mul_out[391][6]);
mul_8x8bit m1175 (image[170],filter[5],mul_out[391][7]);
mul_8x8bit m1176 (image[196],filter[6],mul_out[392][5]);
mul_8x8bit m1177 (image[197],filter[7],mul_out[392][6]);
mul_8x8bit m1178 (image[198],filter[8],mul_out[392][7]);

adder_8bit ad130 (mul_out[390][5],mul_out[390][6],mul_out[390][7],mul_out[391][5],mul_out[391][6],mul_out[391][7],mul_out[392][5],mul_out[392][6],mul_out[392][7],conv_out[130]);



mul_8x8bit m1179 (image[141],filter[0],mul_out[393][5]);
mul_8x8bit m1180 (image[142],filter[1],mul_out[393][6]);
mul_8x8bit m1181 (image[143],filter[2],mul_out[393][7]);
mul_8x8bit m1182 (image[169],filter[3],mul_out[394][5]);
mul_8x8bit m1183 (image[170],filter[4],mul_out[394][6]);
mul_8x8bit m1184 (image[171],filter[5],mul_out[394][7]);
mul_8x8bit m1185 (image[197],filter[6],mul_out[395][5]);
mul_8x8bit m1186 (image[198],filter[7],mul_out[395][6]);
mul_8x8bit m1187 (image[199],filter[8],mul_out[395][7]);

adder_8bit ad131 (mul_out[393][5],mul_out[393][6],mul_out[393][7],mul_out[394][5],mul_out[394][6],mul_out[394][7],mul_out[395][5],mul_out[395][6],mul_out[395][7],conv_out[131]);



mul_8x8bit m1188 (image[142],filter[0],mul_out[396][5]);
mul_8x8bit m1189 (image[143],filter[1],mul_out[396][6]);
mul_8x8bit m1190 (image[144],filter[2],mul_out[396][7]);
mul_8x8bit m1191 (image[170],filter[3],mul_out[397][5]);
mul_8x8bit m1192 (image[171],filter[4],mul_out[397][6]);
mul_8x8bit m1193 (image[172],filter[5],mul_out[397][7]);
mul_8x8bit m1194 (image[198],filter[6],mul_out[398][5]);
mul_8x8bit m1195 (image[199],filter[7],mul_out[398][6]);
mul_8x8bit m1196 (image[200],filter[8],mul_out[398][7]);

adder_8bit ad132 (mul_out[396][5],mul_out[396][6],mul_out[396][7],mul_out[397][5],mul_out[397][6],mul_out[397][7],mul_out[398][5],mul_out[398][6],mul_out[398][7],conv_out[132]);



mul_8x8bit m1197 (image[143],filter[0],mul_out[399][5]);
mul_8x8bit m1198 (image[144],filter[1],mul_out[399][6]);
mul_8x8bit m1199 (image[145],filter[2],mul_out[399][7]);
mul_8x8bit m1200 (image[171],filter[3],mul_out[400][5]);
mul_8x8bit m1201 (image[172],filter[4],mul_out[400][6]);
mul_8x8bit m1202 (image[173],filter[5],mul_out[400][7]);
mul_8x8bit m1203 (image[199],filter[6],mul_out[401][5]);
mul_8x8bit m1204 (image[200],filter[7],mul_out[401][6]);
mul_8x8bit m1205 (image[201],filter[8],mul_out[401][7]);

adder_8bit ad133 (mul_out[399][5],mul_out[399][6],mul_out[399][7],mul_out[400][5],mul_out[400][6],mul_out[400][7],mul_out[401][5],mul_out[401][6],mul_out[401][7],conv_out[133]);



mul_8x8bit m1206 (image[144],filter[0],mul_out[402][5]);
mul_8x8bit m1207 (image[145],filter[1],mul_out[402][6]);
mul_8x8bit m1208 (image[146],filter[2],mul_out[402][7]);
mul_8x8bit m1209 (image[172],filter[3],mul_out[403][5]);
mul_8x8bit m1210 (image[173],filter[4],mul_out[403][6]);
mul_8x8bit m1211 (image[174],filter[5],mul_out[403][7]);
mul_8x8bit m1212 (image[200],filter[6],mul_out[404][5]);
mul_8x8bit m1213 (image[201],filter[7],mul_out[404][6]);
mul_8x8bit m1214 (image[202],filter[8],mul_out[404][7]);

adder_8bit ad134 (mul_out[402][5],mul_out[402][6],mul_out[402][7],mul_out[403][5],mul_out[403][6],mul_out[403][7],mul_out[404][5],mul_out[404][6],mul_out[404][7],conv_out[134]);



mul_8x8bit m1215 (image[145],filter[0],mul_out[405][5]);
mul_8x8bit m1216 (image[146],filter[1],mul_out[405][6]);
mul_8x8bit m1217 (image[147],filter[2],mul_out[405][7]);
mul_8x8bit m1218 (image[173],filter[3],mul_out[406][5]);
mul_8x8bit m1219 (image[174],filter[4],mul_out[406][6]);
mul_8x8bit m1220 (image[175],filter[5],mul_out[406][7]);
mul_8x8bit m1221 (image[201],filter[6],mul_out[407][5]);
mul_8x8bit m1222 (image[202],filter[7],mul_out[407][6]);
mul_8x8bit m1223 (image[203],filter[8],mul_out[407][7]);

adder_8bit ad135 (mul_out[405][5],mul_out[405][6],mul_out[405][7],mul_out[406][5],mul_out[406][6],mul_out[406][7],mul_out[407][5],mul_out[407][6],mul_out[407][7],conv_out[135]);



mul_8x8bit m1224 (image[146],filter[0],mul_out[408][5]);
mul_8x8bit m1225 (image[147],filter[1],mul_out[408][6]);
mul_8x8bit m1226 (image[148],filter[2],mul_out[408][7]);
mul_8x8bit m1227 (image[174],filter[3],mul_out[409][5]);
mul_8x8bit m1228 (image[175],filter[4],mul_out[409][6]);
mul_8x8bit m1229 (image[176],filter[5],mul_out[409][7]);
mul_8x8bit m1230 (image[202],filter[6],mul_out[410][5]);
mul_8x8bit m1231 (image[203],filter[7],mul_out[410][6]);
mul_8x8bit m1232 (image[204],filter[8],mul_out[410][7]);

adder_8bit ad136 (mul_out[408][5],mul_out[408][6],mul_out[408][7],mul_out[409][5],mul_out[409][6],mul_out[409][7],mul_out[410][5],mul_out[410][6],mul_out[410][7],conv_out[136]);



mul_8x8bit m1233 (image[147],filter[0],mul_out[411][5]);
mul_8x8bit m1234 (image[148],filter[1],mul_out[411][6]);
mul_8x8bit m1235 (image[149],filter[2],mul_out[411][7]);
mul_8x8bit m1236 (image[175],filter[3],mul_out[412][5]);
mul_8x8bit m1237 (image[176],filter[4],mul_out[412][6]);
mul_8x8bit m1238 (image[177],filter[5],mul_out[412][7]);
mul_8x8bit m1239 (image[203],filter[6],mul_out[413][5]);
mul_8x8bit m1240 (image[204],filter[7],mul_out[413][6]);
mul_8x8bit m1241 (image[205],filter[8],mul_out[413][7]);

adder_8bit ad137 (mul_out[411][5],mul_out[411][6],mul_out[411][7],mul_out[412][5],mul_out[412][6],mul_out[412][7],mul_out[413][5],mul_out[413][6],mul_out[413][7],conv_out[137]);



mul_8x8bit m1242 (image[148],filter[0],mul_out[414][5]);
mul_8x8bit m1243 (image[149],filter[1],mul_out[414][6]);
mul_8x8bit m1244 (image[150],filter[2],mul_out[414][7]);
mul_8x8bit m1245 (image[176],filter[3],mul_out[415][5]);
mul_8x8bit m1246 (image[177],filter[4],mul_out[415][6]);
mul_8x8bit m1247 (image[178],filter[5],mul_out[415][7]);
mul_8x8bit m1248 (image[204],filter[6],mul_out[416][5]);
mul_8x8bit m1249 (image[205],filter[7],mul_out[416][6]);
mul_8x8bit m1250 (image[206],filter[8],mul_out[416][7]);

adder_8bit ad138 (mul_out[414][5],mul_out[414][6],mul_out[414][7],mul_out[415][5],mul_out[415][6],mul_out[415][7],mul_out[416][5],mul_out[416][6],mul_out[416][7],conv_out[138]);



mul_8x8bit m1251 (image[149],filter[0],mul_out[417][5]);
mul_8x8bit m1252 (image[150],filter[1],mul_out[417][6]);
mul_8x8bit m1253 (image[151],filter[2],mul_out[417][7]);
mul_8x8bit m1254 (image[177],filter[3],mul_out[418][5]);
mul_8x8bit m1255 (image[178],filter[4],mul_out[418][6]);
mul_8x8bit m1256 (image[179],filter[5],mul_out[418][7]);
mul_8x8bit m1257 (image[205],filter[6],mul_out[419][5]);
mul_8x8bit m1258 (image[206],filter[7],mul_out[419][6]);
mul_8x8bit m1259 (image[207],filter[8],mul_out[419][7]);

adder_8bit ad139 (mul_out[417][5],mul_out[417][6],mul_out[417][7],mul_out[418][5],mul_out[418][6],mul_out[418][7],mul_out[419][5],mul_out[419][6],mul_out[419][7],conv_out[139]);



mul_8x8bit m1260 (image[150],filter[0],mul_out[420][5]);
mul_8x8bit m1261 (image[151],filter[1],mul_out[420][6]);
mul_8x8bit m1262 (image[152],filter[2],mul_out[420][7]);
mul_8x8bit m1263 (image[178],filter[3],mul_out[421][5]);
mul_8x8bit m1264 (image[179],filter[4],mul_out[421][6]);
mul_8x8bit m1265 (image[180],filter[5],mul_out[421][7]);
mul_8x8bit m1266 (image[206],filter[6],mul_out[422][5]);
mul_8x8bit m1267 (image[207],filter[7],mul_out[422][6]);
mul_8x8bit m1268 (image[208],filter[8],mul_out[422][7]);

adder_8bit ad140 (mul_out[420][5],mul_out[420][6],mul_out[420][7],mul_out[421][5],mul_out[421][6],mul_out[421][7],mul_out[422][5],mul_out[422][6],mul_out[422][7],conv_out[140]);



mul_8x8bit m1269 (image[151],filter[0],mul_out[423][5]);
mul_8x8bit m1270 (image[152],filter[1],mul_out[423][6]);
mul_8x8bit m1271 (image[153],filter[2],mul_out[423][7]);
mul_8x8bit m1272 (image[179],filter[3],mul_out[424][5]);
mul_8x8bit m1273 (image[180],filter[4],mul_out[424][6]);
mul_8x8bit m1274 (image[181],filter[5],mul_out[424][7]);
mul_8x8bit m1275 (image[207],filter[6],mul_out[425][5]);
mul_8x8bit m1276 (image[208],filter[7],mul_out[425][6]);
mul_8x8bit m1277 (image[209],filter[8],mul_out[425][7]);

adder_8bit ad141 (mul_out[423][5],mul_out[423][6],mul_out[423][7],mul_out[424][5],mul_out[424][6],mul_out[424][7],mul_out[425][5],mul_out[425][6],mul_out[425][7],conv_out[141]);



mul_8x8bit m1278 (image[152],filter[0],mul_out[426][5]);
mul_8x8bit m1279 (image[153],filter[1],mul_out[426][6]);
mul_8x8bit m1280 (image[154],filter[2],mul_out[426][7]);
mul_8x8bit m1281 (image[180],filter[3],mul_out[427][5]);
mul_8x8bit m1282 (image[181],filter[4],mul_out[427][6]);
mul_8x8bit m1283 (image[182],filter[5],mul_out[427][7]);
mul_8x8bit m1284 (image[208],filter[6],mul_out[428][5]);
mul_8x8bit m1285 (image[209],filter[7],mul_out[428][6]);
mul_8x8bit m1286 (image[210],filter[8],mul_out[428][7]);

adder_8bit ad142 (mul_out[426][5],mul_out[426][6],mul_out[426][7],mul_out[427][5],mul_out[427][6],mul_out[427][7],mul_out[428][5],mul_out[428][6],mul_out[428][7],conv_out[142]);



mul_8x8bit m1287 (image[153],filter[0],mul_out[429][5]);
mul_8x8bit m1288 (image[154],filter[1],mul_out[429][6]);
mul_8x8bit m1289 (image[155],filter[2],mul_out[429][7]);
mul_8x8bit m1290 (image[181],filter[3],mul_out[430][5]);
mul_8x8bit m1291 (image[182],filter[4],mul_out[430][6]);
mul_8x8bit m1292 (image[183],filter[5],mul_out[430][7]);
mul_8x8bit m1293 (image[209],filter[6],mul_out[431][5]);
mul_8x8bit m1294 (image[210],filter[7],mul_out[431][6]);
mul_8x8bit m1295 (image[211],filter[8],mul_out[431][7]);

adder_8bit ad143 (mul_out[429][5],mul_out[429][6],mul_out[429][7],mul_out[430][5],mul_out[430][6],mul_out[430][7],mul_out[431][5],mul_out[431][6],mul_out[431][7],conv_out[143]);



mul_8x8bit m1296 (image[154],filter[0],mul_out[432][5]);
mul_8x8bit m1297 (image[155],filter[1],mul_out[432][6]);
mul_8x8bit m1298 (image[156],filter[2],mul_out[432][7]);
mul_8x8bit m1299 (image[182],filter[3],mul_out[433][5]);
mul_8x8bit m1300 (image[183],filter[4],mul_out[433][6]);
mul_8x8bit m1301 (image[184],filter[5],mul_out[433][7]);
mul_8x8bit m1302 (image[210],filter[6],mul_out[434][5]);
mul_8x8bit m1303 (image[211],filter[7],mul_out[434][6]);
mul_8x8bit m1304 (image[212],filter[8],mul_out[434][7]);

adder_8bit ad144 (mul_out[432][5],mul_out[432][6],mul_out[432][7],mul_out[433][5],mul_out[433][6],mul_out[433][7],mul_out[434][5],mul_out[434][6],mul_out[434][7],conv_out[144]);



mul_8x8bit m1305 (image[155],filter[0],mul_out[435][5]);
mul_8x8bit m1306 (image[156],filter[1],mul_out[435][6]);
mul_8x8bit m1307 (image[157],filter[2],mul_out[435][7]);
mul_8x8bit m1308 (image[183],filter[3],mul_out[436][5]);
mul_8x8bit m1309 (image[184],filter[4],mul_out[436][6]);
mul_8x8bit m1310 (image[185],filter[5],mul_out[436][7]);
mul_8x8bit m1311 (image[211],filter[6],mul_out[437][5]);
mul_8x8bit m1312 (image[212],filter[7],mul_out[437][6]);
mul_8x8bit m1313 (image[213],filter[8],mul_out[437][7]);

adder_8bit ad145 (mul_out[435][5],mul_out[435][6],mul_out[435][7],mul_out[436][5],mul_out[436][6],mul_out[436][7],mul_out[437][5],mul_out[437][6],mul_out[437][7],conv_out[145]);



mul_8x8bit m1314 (image[156],filter[0],mul_out[438][5]);
mul_8x8bit m1315 (image[157],filter[1],mul_out[438][6]);
mul_8x8bit m1316 (image[158],filter[2],mul_out[438][7]);
mul_8x8bit m1317 (image[184],filter[3],mul_out[439][5]);
mul_8x8bit m1318 (image[185],filter[4],mul_out[439][6]);
mul_8x8bit m1319 (image[186],filter[5],mul_out[439][7]);
mul_8x8bit m1320 (image[212],filter[6],mul_out[440][5]);
mul_8x8bit m1321 (image[213],filter[7],mul_out[440][6]);
mul_8x8bit m1322 (image[214],filter[8],mul_out[440][7]);

adder_8bit ad146 (mul_out[438][5],mul_out[438][6],mul_out[438][7],mul_out[439][5],mul_out[439][6],mul_out[439][7],mul_out[440][5],mul_out[440][6],mul_out[440][7],conv_out[146]);



mul_8x8bit m1323 (image[157],filter[0],mul_out[441][5]);
mul_8x8bit m1324 (image[158],filter[1],mul_out[441][6]);
mul_8x8bit m1325 (image[159],filter[2],mul_out[441][7]);
mul_8x8bit m1326 (image[185],filter[3],mul_out[442][5]);
mul_8x8bit m1327 (image[186],filter[4],mul_out[442][6]);
mul_8x8bit m1328 (image[187],filter[5],mul_out[442][7]);
mul_8x8bit m1329 (image[213],filter[6],mul_out[443][5]);
mul_8x8bit m1330 (image[214],filter[7],mul_out[443][6]);
mul_8x8bit m1331 (image[215],filter[8],mul_out[443][7]);

adder_8bit ad147 (mul_out[441][5],mul_out[441][6],mul_out[441][7],mul_out[442][5],mul_out[442][6],mul_out[442][7],mul_out[443][5],mul_out[443][6],mul_out[443][7],conv_out[147]);



mul_8x8bit m1332 (image[158],filter[0],mul_out[444][5]);
mul_8x8bit m1333 (image[159],filter[1],mul_out[444][6]);
mul_8x8bit m1334 (image[160],filter[2],mul_out[444][7]);
mul_8x8bit m1335 (image[186],filter[3],mul_out[445][5]);
mul_8x8bit m1336 (image[187],filter[4],mul_out[445][6]);
mul_8x8bit m1337 (image[188],filter[5],mul_out[445][7]);
mul_8x8bit m1338 (image[214],filter[6],mul_out[446][5]);
mul_8x8bit m1339 (image[215],filter[7],mul_out[446][6]);
mul_8x8bit m1340 (image[216],filter[8],mul_out[446][7]);

adder_8bit ad148 (mul_out[444][5],mul_out[444][6],mul_out[444][7],mul_out[445][5],mul_out[445][6],mul_out[445][7],mul_out[446][5],mul_out[446][6],mul_out[446][7],conv_out[148]);



mul_8x8bit m1341 (image[159],filter[0],mul_out[447][5]);
mul_8x8bit m1342 (image[160],filter[1],mul_out[447][6]);
mul_8x8bit m1343 (image[161],filter[2],mul_out[447][7]);
mul_8x8bit m1344 (image[187],filter[3],mul_out[448][5]);
mul_8x8bit m1345 (image[188],filter[4],mul_out[448][6]);
mul_8x8bit m1346 (image[189],filter[5],mul_out[448][7]);
mul_8x8bit m1347 (image[215],filter[6],mul_out[449][5]);
mul_8x8bit m1348 (image[216],filter[7],mul_out[449][6]);
mul_8x8bit m1349 (image[217],filter[8],mul_out[449][7]);

adder_8bit ad149 (mul_out[447][5],mul_out[447][6],mul_out[447][7],mul_out[448][5],mul_out[448][6],mul_out[448][7],mul_out[449][5],mul_out[449][6],mul_out[449][7],conv_out[149]);



mul_8x8bit m1350 (image[160],filter[0],mul_out[450][5]);
mul_8x8bit m1351 (image[161],filter[1],mul_out[450][6]);
mul_8x8bit m1352 (image[162],filter[2],mul_out[450][7]);
mul_8x8bit m1353 (image[188],filter[3],mul_out[451][5]);
mul_8x8bit m1354 (image[189],filter[4],mul_out[451][6]);
mul_8x8bit m1355 (image[190],filter[5],mul_out[451][7]);
mul_8x8bit m1356 (image[216],filter[6],mul_out[452][5]);
mul_8x8bit m1357 (image[217],filter[7],mul_out[452][6]);
mul_8x8bit m1358 (image[218],filter[8],mul_out[452][7]);

adder_8bit ad150 (mul_out[450][5],mul_out[450][6],mul_out[450][7],mul_out[451][5],mul_out[451][6],mul_out[451][7],mul_out[452][5],mul_out[452][6],mul_out[452][7],conv_out[150]);



mul_8x8bit m1359 (image[161],filter[0],mul_out[453][5]);
mul_8x8bit m1360 (image[162],filter[1],mul_out[453][6]);
mul_8x8bit m1361 (image[163],filter[2],mul_out[453][7]);
mul_8x8bit m1362 (image[189],filter[3],mul_out[454][5]);
mul_8x8bit m1363 (image[190],filter[4],mul_out[454][6]);
mul_8x8bit m1364 (image[191],filter[5],mul_out[454][7]);
mul_8x8bit m1365 (image[217],filter[6],mul_out[455][5]);
mul_8x8bit m1366 (image[218],filter[7],mul_out[455][6]);
mul_8x8bit m1367 (image[219],filter[8],mul_out[455][7]);

adder_8bit ad151 (mul_out[453][5],mul_out[453][6],mul_out[453][7],mul_out[454][5],mul_out[454][6],mul_out[454][7],mul_out[455][5],mul_out[455][6],mul_out[455][7],conv_out[151]);



mul_8x8bit m1368 (image[162],filter[0],mul_out[456][5]);
mul_8x8bit m1369 (image[163],filter[1],mul_out[456][6]);
mul_8x8bit m1370 (image[164],filter[2],mul_out[456][7]);
mul_8x8bit m1371 (image[190],filter[3],mul_out[457][5]);
mul_8x8bit m1372 (image[191],filter[4],mul_out[457][6]);
mul_8x8bit m1373 (image[192],filter[5],mul_out[457][7]);
mul_8x8bit m1374 (image[218],filter[6],mul_out[458][5]);
mul_8x8bit m1375 (image[219],filter[7],mul_out[458][6]);
mul_8x8bit m1376 (image[220],filter[8],mul_out[458][7]);

adder_8bit ad152 (mul_out[456][5],mul_out[456][6],mul_out[456][7],mul_out[457][5],mul_out[457][6],mul_out[457][7],mul_out[458][5],mul_out[458][6],mul_out[458][7],conv_out[152]);



mul_8x8bit m1377 (image[163],filter[0],mul_out[459][5]);
mul_8x8bit m1378 (image[164],filter[1],mul_out[459][6]);
mul_8x8bit m1379 (image[165],filter[2],mul_out[459][7]);
mul_8x8bit m1380 (image[191],filter[3],mul_out[460][5]);
mul_8x8bit m1381 (image[192],filter[4],mul_out[460][6]);
mul_8x8bit m1382 (image[193],filter[5],mul_out[460][7]);
mul_8x8bit m1383 (image[219],filter[6],mul_out[461][5]);
mul_8x8bit m1384 (image[220],filter[7],mul_out[461][6]);
mul_8x8bit m1385 (image[221],filter[8],mul_out[461][7]);

adder_8bit ad153 (mul_out[459][5],mul_out[459][6],mul_out[459][7],mul_out[460][5],mul_out[460][6],mul_out[460][7],mul_out[461][5],mul_out[461][6],mul_out[461][7],conv_out[153]);



mul_8x8bit m1386 (image[164],filter[0],mul_out[462][5]);
mul_8x8bit m1387 (image[165],filter[1],mul_out[462][6]);
mul_8x8bit m1388 (image[166],filter[2],mul_out[462][7]);
mul_8x8bit m1389 (image[192],filter[3],mul_out[463][5]);
mul_8x8bit m1390 (image[193],filter[4],mul_out[463][6]);
mul_8x8bit m1391 (image[194],filter[5],mul_out[463][7]);
mul_8x8bit m1392 (image[220],filter[6],mul_out[464][5]);
mul_8x8bit m1393 (image[221],filter[7],mul_out[464][6]);
mul_8x8bit m1394 (image[222],filter[8],mul_out[464][7]);

adder_8bit ad154 (mul_out[462][5],mul_out[462][6],mul_out[462][7],mul_out[463][5],mul_out[463][6],mul_out[463][7],mul_out[464][5],mul_out[464][6],mul_out[464][7],conv_out[154]);



mul_8x8bit m1395 (image[165],filter[0],mul_out[465][5]);
mul_8x8bit m1396 (image[166],filter[1],mul_out[465][6]);
mul_8x8bit m1397 (image[167],filter[2],mul_out[465][7]);
mul_8x8bit m1398 (image[193],filter[3],mul_out[466][5]);
mul_8x8bit m1399 (image[194],filter[4],mul_out[466][6]);
mul_8x8bit m1400 (image[195],filter[5],mul_out[466][7]);
mul_8x8bit m1401 (image[221],filter[6],mul_out[467][5]);
mul_8x8bit m1402 (image[222],filter[7],mul_out[467][6]);
mul_8x8bit m1403 (image[223],filter[8],mul_out[467][7]);

adder_8bit ad155 (mul_out[465][5],mul_out[465][6],mul_out[465][7],mul_out[466][5],mul_out[466][6],mul_out[466][7],mul_out[467][5],mul_out[467][6],mul_out[467][7],conv_out[155]);



mul_8x8bit m1404 (image[168],filter[0],mul_out[468][6]);
mul_8x8bit m1405 (image[169],filter[1],mul_out[468][7]);
mul_8x8bit m1406 (image[170],filter[2],mul_out[468][8]);
mul_8x8bit m1407 (image[196],filter[3],mul_out[469][6]);
mul_8x8bit m1408 (image[197],filter[4],mul_out[469][7]);
mul_8x8bit m1409 (image[198],filter[5],mul_out[469][8]);
mul_8x8bit m1410 (image[224],filter[6],mul_out[470][6]);
mul_8x8bit m1411 (image[225],filter[7],mul_out[470][7]);
mul_8x8bit m1412 (image[226],filter[8],mul_out[470][8]);

adder_8bit ad156 (mul_out[468][6],mul_out[468][7],mul_out[468][8],mul_out[469][6],mul_out[469][7],mul_out[469][8],mul_out[470][6],mul_out[470][7],mul_out[470][8],conv_out[156]);



mul_8x8bit m1413 (image[169],filter[0],mul_out[471][6]);
mul_8x8bit m1414 (image[170],filter[1],mul_out[471][7]);
mul_8x8bit m1415 (image[171],filter[2],mul_out[471][8]);
mul_8x8bit m1416 (image[197],filter[3],mul_out[472][6]);
mul_8x8bit m1417 (image[198],filter[4],mul_out[472][7]);
mul_8x8bit m1418 (image[199],filter[5],mul_out[472][8]);
mul_8x8bit m1419 (image[225],filter[6],mul_out[473][6]);
mul_8x8bit m1420 (image[226],filter[7],mul_out[473][7]);
mul_8x8bit m1421 (image[227],filter[8],mul_out[473][8]);

adder_8bit ad157 (mul_out[471][6],mul_out[471][7],mul_out[471][8],mul_out[472][6],mul_out[472][7],mul_out[472][8],mul_out[473][6],mul_out[473][7],mul_out[473][8],conv_out[157]);



mul_8x8bit m1422 (image[170],filter[0],mul_out[474][6]);
mul_8x8bit m1423 (image[171],filter[1],mul_out[474][7]);
mul_8x8bit m1424 (image[172],filter[2],mul_out[474][8]);
mul_8x8bit m1425 (image[198],filter[3],mul_out[475][6]);
mul_8x8bit m1426 (image[199],filter[4],mul_out[475][7]);
mul_8x8bit m1427 (image[200],filter[5],mul_out[475][8]);
mul_8x8bit m1428 (image[226],filter[6],mul_out[476][6]);
mul_8x8bit m1429 (image[227],filter[7],mul_out[476][7]);
mul_8x8bit m1430 (image[228],filter[8],mul_out[476][8]);

adder_8bit ad158 (mul_out[474][6],mul_out[474][7],mul_out[474][8],mul_out[475][6],mul_out[475][7],mul_out[475][8],mul_out[476][6],mul_out[476][7],mul_out[476][8],conv_out[158]);



mul_8x8bit m1431 (image[171],filter[0],mul_out[477][6]);
mul_8x8bit m1432 (image[172],filter[1],mul_out[477][7]);
mul_8x8bit m1433 (image[173],filter[2],mul_out[477][8]);
mul_8x8bit m1434 (image[199],filter[3],mul_out[478][6]);
mul_8x8bit m1435 (image[200],filter[4],mul_out[478][7]);
mul_8x8bit m1436 (image[201],filter[5],mul_out[478][8]);
mul_8x8bit m1437 (image[227],filter[6],mul_out[479][6]);
mul_8x8bit m1438 (image[228],filter[7],mul_out[479][7]);
mul_8x8bit m1439 (image[229],filter[8],mul_out[479][8]);

adder_8bit ad159 (mul_out[477][6],mul_out[477][7],mul_out[477][8],mul_out[478][6],mul_out[478][7],mul_out[478][8],mul_out[479][6],mul_out[479][7],mul_out[479][8],conv_out[159]);



mul_8x8bit m1440 (image[172],filter[0],mul_out[480][6]);
mul_8x8bit m1441 (image[173],filter[1],mul_out[480][7]);
mul_8x8bit m1442 (image[174],filter[2],mul_out[480][8]);
mul_8x8bit m1443 (image[200],filter[3],mul_out[481][6]);
mul_8x8bit m1444 (image[201],filter[4],mul_out[481][7]);
mul_8x8bit m1445 (image[202],filter[5],mul_out[481][8]);
mul_8x8bit m1446 (image[228],filter[6],mul_out[482][6]);
mul_8x8bit m1447 (image[229],filter[7],mul_out[482][7]);
mul_8x8bit m1448 (image[230],filter[8],mul_out[482][8]);

adder_8bit ad160 (mul_out[480][6],mul_out[480][7],mul_out[480][8],mul_out[481][6],mul_out[481][7],mul_out[481][8],mul_out[482][6],mul_out[482][7],mul_out[482][8],conv_out[160]);



mul_8x8bit m1449 (image[173],filter[0],mul_out[483][6]);
mul_8x8bit m1450 (image[174],filter[1],mul_out[483][7]);
mul_8x8bit m1451 (image[175],filter[2],mul_out[483][8]);
mul_8x8bit m1452 (image[201],filter[3],mul_out[484][6]);
mul_8x8bit m1453 (image[202],filter[4],mul_out[484][7]);
mul_8x8bit m1454 (image[203],filter[5],mul_out[484][8]);
mul_8x8bit m1455 (image[229],filter[6],mul_out[485][6]);
mul_8x8bit m1456 (image[230],filter[7],mul_out[485][7]);
mul_8x8bit m1457 (image[231],filter[8],mul_out[485][8]);

adder_8bit ad161 (mul_out[483][6],mul_out[483][7],mul_out[483][8],mul_out[484][6],mul_out[484][7],mul_out[484][8],mul_out[485][6],mul_out[485][7],mul_out[485][8],conv_out[161]);



mul_8x8bit m1458 (image[174],filter[0],mul_out[486][6]);
mul_8x8bit m1459 (image[175],filter[1],mul_out[486][7]);
mul_8x8bit m1460 (image[176],filter[2],mul_out[486][8]);
mul_8x8bit m1461 (image[202],filter[3],mul_out[487][6]);
mul_8x8bit m1462 (image[203],filter[4],mul_out[487][7]);
mul_8x8bit m1463 (image[204],filter[5],mul_out[487][8]);
mul_8x8bit m1464 (image[230],filter[6],mul_out[488][6]);
mul_8x8bit m1465 (image[231],filter[7],mul_out[488][7]);
mul_8x8bit m1466 (image[232],filter[8],mul_out[488][8]);

adder_8bit ad162 (mul_out[486][6],mul_out[486][7],mul_out[486][8],mul_out[487][6],mul_out[487][7],mul_out[487][8],mul_out[488][6],mul_out[488][7],mul_out[488][8],conv_out[162]);



mul_8x8bit m1467 (image[175],filter[0],mul_out[489][6]);
mul_8x8bit m1468 (image[176],filter[1],mul_out[489][7]);
mul_8x8bit m1469 (image[177],filter[2],mul_out[489][8]);
mul_8x8bit m1470 (image[203],filter[3],mul_out[490][6]);
mul_8x8bit m1471 (image[204],filter[4],mul_out[490][7]);
mul_8x8bit m1472 (image[205],filter[5],mul_out[490][8]);
mul_8x8bit m1473 (image[231],filter[6],mul_out[491][6]);
mul_8x8bit m1474 (image[232],filter[7],mul_out[491][7]);
mul_8x8bit m1475 (image[233],filter[8],mul_out[491][8]);

adder_8bit ad163 (mul_out[489][6],mul_out[489][7],mul_out[489][8],mul_out[490][6],mul_out[490][7],mul_out[490][8],mul_out[491][6],mul_out[491][7],mul_out[491][8],conv_out[163]);



mul_8x8bit m1476 (image[176],filter[0],mul_out[492][6]);
mul_8x8bit m1477 (image[177],filter[1],mul_out[492][7]);
mul_8x8bit m1478 (image[178],filter[2],mul_out[492][8]);
mul_8x8bit m1479 (image[204],filter[3],mul_out[493][6]);
mul_8x8bit m1480 (image[205],filter[4],mul_out[493][7]);
mul_8x8bit m1481 (image[206],filter[5],mul_out[493][8]);
mul_8x8bit m1482 (image[232],filter[6],mul_out[494][6]);
mul_8x8bit m1483 (image[233],filter[7],mul_out[494][7]);
mul_8x8bit m1484 (image[234],filter[8],mul_out[494][8]);

adder_8bit ad164 (mul_out[492][6],mul_out[492][7],mul_out[492][8],mul_out[493][6],mul_out[493][7],mul_out[493][8],mul_out[494][6],mul_out[494][7],mul_out[494][8],conv_out[164]);



mul_8x8bit m1485 (image[177],filter[0],mul_out[495][6]);
mul_8x8bit m1486 (image[178],filter[1],mul_out[495][7]);
mul_8x8bit m1487 (image[179],filter[2],mul_out[495][8]);
mul_8x8bit m1488 (image[205],filter[3],mul_out[496][6]);
mul_8x8bit m1489 (image[206],filter[4],mul_out[496][7]);
mul_8x8bit m1490 (image[207],filter[5],mul_out[496][8]);
mul_8x8bit m1491 (image[233],filter[6],mul_out[497][6]);
mul_8x8bit m1492 (image[234],filter[7],mul_out[497][7]);
mul_8x8bit m1493 (image[235],filter[8],mul_out[497][8]);

adder_8bit ad165 (mul_out[495][6],mul_out[495][7],mul_out[495][8],mul_out[496][6],mul_out[496][7],mul_out[496][8],mul_out[497][6],mul_out[497][7],mul_out[497][8],conv_out[165]);



mul_8x8bit m1494 (image[178],filter[0],mul_out[498][6]);
mul_8x8bit m1495 (image[179],filter[1],mul_out[498][7]);
mul_8x8bit m1496 (image[180],filter[2],mul_out[498][8]);
mul_8x8bit m1497 (image[206],filter[3],mul_out[499][6]);
mul_8x8bit m1498 (image[207],filter[4],mul_out[499][7]);
mul_8x8bit m1499 (image[208],filter[5],mul_out[499][8]);
mul_8x8bit m1500 (image[234],filter[6],mul_out[500][6]);
mul_8x8bit m1501 (image[235],filter[7],mul_out[500][7]);
mul_8x8bit m1502 (image[236],filter[8],mul_out[500][8]);

adder_8bit ad166 (mul_out[498][6],mul_out[498][7],mul_out[498][8],mul_out[499][6],mul_out[499][7],mul_out[499][8],mul_out[500][6],mul_out[500][7],mul_out[500][8],conv_out[166]);



mul_8x8bit m1503 (image[179],filter[0],mul_out[501][6]);
mul_8x8bit m1504 (image[180],filter[1],mul_out[501][7]);
mul_8x8bit m1505 (image[181],filter[2],mul_out[501][8]);
mul_8x8bit m1506 (image[207],filter[3],mul_out[502][6]);
mul_8x8bit m1507 (image[208],filter[4],mul_out[502][7]);
mul_8x8bit m1508 (image[209],filter[5],mul_out[502][8]);
mul_8x8bit m1509 (image[235],filter[6],mul_out[503][6]);
mul_8x8bit m1510 (image[236],filter[7],mul_out[503][7]);
mul_8x8bit m1511 (image[237],filter[8],mul_out[503][8]);

adder_8bit ad167 (mul_out[501][6],mul_out[501][7],mul_out[501][8],mul_out[502][6],mul_out[502][7],mul_out[502][8],mul_out[503][6],mul_out[503][7],mul_out[503][8],conv_out[167]);



mul_8x8bit m1512 (image[180],filter[0],mul_out[504][6]);
mul_8x8bit m1513 (image[181],filter[1],mul_out[504][7]);
mul_8x8bit m1514 (image[182],filter[2],mul_out[504][8]);
mul_8x8bit m1515 (image[208],filter[3],mul_out[505][6]);
mul_8x8bit m1516 (image[209],filter[4],mul_out[505][7]);
mul_8x8bit m1517 (image[210],filter[5],mul_out[505][8]);
mul_8x8bit m1518 (image[236],filter[6],mul_out[506][6]);
mul_8x8bit m1519 (image[237],filter[7],mul_out[506][7]);
mul_8x8bit m1520 (image[238],filter[8],mul_out[506][8]);

adder_8bit ad168 (mul_out[504][6],mul_out[504][7],mul_out[504][8],mul_out[505][6],mul_out[505][7],mul_out[505][8],mul_out[506][6],mul_out[506][7],mul_out[506][8],conv_out[168]);



mul_8x8bit m1521 (image[181],filter[0],mul_out[507][6]);
mul_8x8bit m1522 (image[182],filter[1],mul_out[507][7]);
mul_8x8bit m1523 (image[183],filter[2],mul_out[507][8]);
mul_8x8bit m1524 (image[209],filter[3],mul_out[508][6]);
mul_8x8bit m1525 (image[210],filter[4],mul_out[508][7]);
mul_8x8bit m1526 (image[211],filter[5],mul_out[508][8]);
mul_8x8bit m1527 (image[237],filter[6],mul_out[509][6]);
mul_8x8bit m1528 (image[238],filter[7],mul_out[509][7]);
mul_8x8bit m1529 (image[239],filter[8],mul_out[509][8]);

adder_8bit ad169 (mul_out[507][6],mul_out[507][7],mul_out[507][8],mul_out[508][6],mul_out[508][7],mul_out[508][8],mul_out[509][6],mul_out[509][7],mul_out[509][8],conv_out[169]);



mul_8x8bit m1530 (image[182],filter[0],mul_out[510][6]);
mul_8x8bit m1531 (image[183],filter[1],mul_out[510][7]);
mul_8x8bit m1532 (image[184],filter[2],mul_out[510][8]);
mul_8x8bit m1533 (image[210],filter[3],mul_out[511][6]);
mul_8x8bit m1534 (image[211],filter[4],mul_out[511][7]);
mul_8x8bit m1535 (image[212],filter[5],mul_out[511][8]);
mul_8x8bit m1536 (image[238],filter[6],mul_out[512][6]);
mul_8x8bit m1537 (image[239],filter[7],mul_out[512][7]);
mul_8x8bit m1538 (image[240],filter[8],mul_out[512][8]);

adder_8bit ad170 (mul_out[510][6],mul_out[510][7],mul_out[510][8],mul_out[511][6],mul_out[511][7],mul_out[511][8],mul_out[512][6],mul_out[512][7],mul_out[512][8],conv_out[170]);



mul_8x8bit m1539 (image[183],filter[0],mul_out[513][6]);
mul_8x8bit m1540 (image[184],filter[1],mul_out[513][7]);
mul_8x8bit m1541 (image[185],filter[2],mul_out[513][8]);
mul_8x8bit m1542 (image[211],filter[3],mul_out[514][6]);
mul_8x8bit m1543 (image[212],filter[4],mul_out[514][7]);
mul_8x8bit m1544 (image[213],filter[5],mul_out[514][8]);
mul_8x8bit m1545 (image[239],filter[6],mul_out[515][6]);
mul_8x8bit m1546 (image[240],filter[7],mul_out[515][7]);
mul_8x8bit m1547 (image[241],filter[8],mul_out[515][8]);

adder_8bit ad171 (mul_out[513][6],mul_out[513][7],mul_out[513][8],mul_out[514][6],mul_out[514][7],mul_out[514][8],mul_out[515][6],mul_out[515][7],mul_out[515][8],conv_out[171]);



mul_8x8bit m1548 (image[184],filter[0],mul_out[516][6]);
mul_8x8bit m1549 (image[185],filter[1],mul_out[516][7]);
mul_8x8bit m1550 (image[186],filter[2],mul_out[516][8]);
mul_8x8bit m1551 (image[212],filter[3],mul_out[517][6]);
mul_8x8bit m1552 (image[213],filter[4],mul_out[517][7]);
mul_8x8bit m1553 (image[214],filter[5],mul_out[517][8]);
mul_8x8bit m1554 (image[240],filter[6],mul_out[518][6]);
mul_8x8bit m1555 (image[241],filter[7],mul_out[518][7]);
mul_8x8bit m1556 (image[242],filter[8],mul_out[518][8]);

adder_8bit ad172 (mul_out[516][6],mul_out[516][7],mul_out[516][8],mul_out[517][6],mul_out[517][7],mul_out[517][8],mul_out[518][6],mul_out[518][7],mul_out[518][8],conv_out[172]);



mul_8x8bit m1557 (image[185],filter[0],mul_out[519][6]);
mul_8x8bit m1558 (image[186],filter[1],mul_out[519][7]);
mul_8x8bit m1559 (image[187],filter[2],mul_out[519][8]);
mul_8x8bit m1560 (image[213],filter[3],mul_out[520][6]);
mul_8x8bit m1561 (image[214],filter[4],mul_out[520][7]);
mul_8x8bit m1562 (image[215],filter[5],mul_out[520][8]);
mul_8x8bit m1563 (image[241],filter[6],mul_out[521][6]);
mul_8x8bit m1564 (image[242],filter[7],mul_out[521][7]);
mul_8x8bit m1565 (image[243],filter[8],mul_out[521][8]);

adder_8bit ad173 (mul_out[519][6],mul_out[519][7],mul_out[519][8],mul_out[520][6],mul_out[520][7],mul_out[520][8],mul_out[521][6],mul_out[521][7],mul_out[521][8],conv_out[173]);



mul_8x8bit m1566 (image[186],filter[0],mul_out[522][6]);
mul_8x8bit m1567 (image[187],filter[1],mul_out[522][7]);
mul_8x8bit m1568 (image[188],filter[2],mul_out[522][8]);
mul_8x8bit m1569 (image[214],filter[3],mul_out[523][6]);
mul_8x8bit m1570 (image[215],filter[4],mul_out[523][7]);
mul_8x8bit m1571 (image[216],filter[5],mul_out[523][8]);
mul_8x8bit m1572 (image[242],filter[6],mul_out[524][6]);
mul_8x8bit m1573 (image[243],filter[7],mul_out[524][7]);
mul_8x8bit m1574 (image[244],filter[8],mul_out[524][8]);

adder_8bit ad174 (mul_out[522][6],mul_out[522][7],mul_out[522][8],mul_out[523][6],mul_out[523][7],mul_out[523][8],mul_out[524][6],mul_out[524][7],mul_out[524][8],conv_out[174]);



mul_8x8bit m1575 (image[187],filter[0],mul_out[525][6]);
mul_8x8bit m1576 (image[188],filter[1],mul_out[525][7]);
mul_8x8bit m1577 (image[189],filter[2],mul_out[525][8]);
mul_8x8bit m1578 (image[215],filter[3],mul_out[526][6]);
mul_8x8bit m1579 (image[216],filter[4],mul_out[526][7]);
mul_8x8bit m1580 (image[217],filter[5],mul_out[526][8]);
mul_8x8bit m1581 (image[243],filter[6],mul_out[527][6]);
mul_8x8bit m1582 (image[244],filter[7],mul_out[527][7]);
mul_8x8bit m1583 (image[245],filter[8],mul_out[527][8]);

adder_8bit ad175 (mul_out[525][6],mul_out[525][7],mul_out[525][8],mul_out[526][6],mul_out[526][7],mul_out[526][8],mul_out[527][6],mul_out[527][7],mul_out[527][8],conv_out[175]);



mul_8x8bit m1584 (image[188],filter[0],mul_out[528][6]);
mul_8x8bit m1585 (image[189],filter[1],mul_out[528][7]);
mul_8x8bit m1586 (image[190],filter[2],mul_out[528][8]);
mul_8x8bit m1587 (image[216],filter[3],mul_out[529][6]);
mul_8x8bit m1588 (image[217],filter[4],mul_out[529][7]);
mul_8x8bit m1589 (image[218],filter[5],mul_out[529][8]);
mul_8x8bit m1590 (image[244],filter[6],mul_out[530][6]);
mul_8x8bit m1591 (image[245],filter[7],mul_out[530][7]);
mul_8x8bit m1592 (image[246],filter[8],mul_out[530][8]);

adder_8bit ad176 (mul_out[528][6],mul_out[528][7],mul_out[528][8],mul_out[529][6],mul_out[529][7],mul_out[529][8],mul_out[530][6],mul_out[530][7],mul_out[530][8],conv_out[176]);



mul_8x8bit m1593 (image[189],filter[0],mul_out[531][6]);
mul_8x8bit m1594 (image[190],filter[1],mul_out[531][7]);
mul_8x8bit m1595 (image[191],filter[2],mul_out[531][8]);
mul_8x8bit m1596 (image[217],filter[3],mul_out[532][6]);
mul_8x8bit m1597 (image[218],filter[4],mul_out[532][7]);
mul_8x8bit m1598 (image[219],filter[5],mul_out[532][8]);
mul_8x8bit m1599 (image[245],filter[6],mul_out[533][6]);
mul_8x8bit m1600 (image[246],filter[7],mul_out[533][7]);
mul_8x8bit m1601 (image[247],filter[8],mul_out[533][8]);

adder_8bit ad177 (mul_out[531][6],mul_out[531][7],mul_out[531][8],mul_out[532][6],mul_out[532][7],mul_out[532][8],mul_out[533][6],mul_out[533][7],mul_out[533][8],conv_out[177]);



mul_8x8bit m1602 (image[190],filter[0],mul_out[534][6]);
mul_8x8bit m1603 (image[191],filter[1],mul_out[534][7]);
mul_8x8bit m1604 (image[192],filter[2],mul_out[534][8]);
mul_8x8bit m1605 (image[218],filter[3],mul_out[535][6]);
mul_8x8bit m1606 (image[219],filter[4],mul_out[535][7]);
mul_8x8bit m1607 (image[220],filter[5],mul_out[535][8]);
mul_8x8bit m1608 (image[246],filter[6],mul_out[536][6]);
mul_8x8bit m1609 (image[247],filter[7],mul_out[536][7]);
mul_8x8bit m1610 (image[248],filter[8],mul_out[536][8]);

adder_8bit ad178 (mul_out[534][6],mul_out[534][7],mul_out[534][8],mul_out[535][6],mul_out[535][7],mul_out[535][8],mul_out[536][6],mul_out[536][7],mul_out[536][8],conv_out[178]);



mul_8x8bit m1611 (image[191],filter[0],mul_out[537][6]);
mul_8x8bit m1612 (image[192],filter[1],mul_out[537][7]);
mul_8x8bit m1613 (image[193],filter[2],mul_out[537][8]);
mul_8x8bit m1614 (image[219],filter[3],mul_out[538][6]);
mul_8x8bit m1615 (image[220],filter[4],mul_out[538][7]);
mul_8x8bit m1616 (image[221],filter[5],mul_out[538][8]);
mul_8x8bit m1617 (image[247],filter[6],mul_out[539][6]);
mul_8x8bit m1618 (image[248],filter[7],mul_out[539][7]);
mul_8x8bit m1619 (image[249],filter[8],mul_out[539][8]);

adder_8bit ad179 (mul_out[537][6],mul_out[537][7],mul_out[537][8],mul_out[538][6],mul_out[538][7],mul_out[538][8],mul_out[539][6],mul_out[539][7],mul_out[539][8],conv_out[179]);



mul_8x8bit m1620 (image[192],filter[0],mul_out[540][6]);
mul_8x8bit m1621 (image[193],filter[1],mul_out[540][7]);
mul_8x8bit m1622 (image[194],filter[2],mul_out[540][8]);
mul_8x8bit m1623 (image[220],filter[3],mul_out[541][6]);
mul_8x8bit m1624 (image[221],filter[4],mul_out[541][7]);
mul_8x8bit m1625 (image[222],filter[5],mul_out[541][8]);
mul_8x8bit m1626 (image[248],filter[6],mul_out[542][6]);
mul_8x8bit m1627 (image[249],filter[7],mul_out[542][7]);
mul_8x8bit m1628 (image[250],filter[8],mul_out[542][8]);

adder_8bit ad180 (mul_out[540][6],mul_out[540][7],mul_out[540][8],mul_out[541][6],mul_out[541][7],mul_out[541][8],mul_out[542][6],mul_out[542][7],mul_out[542][8],conv_out[180]);



mul_8x8bit m1629 (image[193],filter[0],mul_out[543][6]);
mul_8x8bit m1630 (image[194],filter[1],mul_out[543][7]);
mul_8x8bit m1631 (image[195],filter[2],mul_out[543][8]);
mul_8x8bit m1632 (image[221],filter[3],mul_out[544][6]);
mul_8x8bit m1633 (image[222],filter[4],mul_out[544][7]);
mul_8x8bit m1634 (image[223],filter[5],mul_out[544][8]);
mul_8x8bit m1635 (image[249],filter[6],mul_out[545][6]);
mul_8x8bit m1636 (image[250],filter[7],mul_out[545][7]);
mul_8x8bit m1637 (image[251],filter[8],mul_out[545][8]);

adder_8bit ad181 (mul_out[543][6],mul_out[543][7],mul_out[543][8],mul_out[544][6],mul_out[544][7],mul_out[544][8],mul_out[545][6],mul_out[545][7],mul_out[545][8],conv_out[181]);



mul_8x8bit m1638 (image[196],filter[0],mul_out[546][7]);
mul_8x8bit m1639 (image[197],filter[1],mul_out[546][8]);
mul_8x8bit m1640 (image[198],filter[2],mul_out[546][9]);
mul_8x8bit m1641 (image[224],filter[3],mul_out[547][7]);
mul_8x8bit m1642 (image[225],filter[4],mul_out[547][8]);
mul_8x8bit m1643 (image[226],filter[5],mul_out[547][9]);
mul_8x8bit m1644 (image[252],filter[6],mul_out[548][7]);
mul_8x8bit m1645 (image[253],filter[7],mul_out[548][8]);
mul_8x8bit m1646 (image[254],filter[8],mul_out[548][9]);

adder_8bit ad182 (mul_out[546][7],mul_out[546][8],mul_out[546][9],mul_out[547][7],mul_out[547][8],mul_out[547][9],mul_out[548][7],mul_out[548][8],mul_out[548][9],conv_out[182]);



mul_8x8bit m1647 (image[197],filter[0],mul_out[549][7]);
mul_8x8bit m1648 (image[198],filter[1],mul_out[549][8]);
mul_8x8bit m1649 (image[199],filter[2],mul_out[549][9]);
mul_8x8bit m1650 (image[225],filter[3],mul_out[550][7]);
mul_8x8bit m1651 (image[226],filter[4],mul_out[550][8]);
mul_8x8bit m1652 (image[227],filter[5],mul_out[550][9]);
mul_8x8bit m1653 (image[253],filter[6],mul_out[551][7]);
mul_8x8bit m1654 (image[254],filter[7],mul_out[551][8]);
mul_8x8bit m1655 (image[255],filter[8],mul_out[551][9]);

adder_8bit ad183 (mul_out[549][7],mul_out[549][8],mul_out[549][9],mul_out[550][7],mul_out[550][8],mul_out[550][9],mul_out[551][7],mul_out[551][8],mul_out[551][9],conv_out[183]);



mul_8x8bit m1656 (image[198],filter[0],mul_out[552][7]);
mul_8x8bit m1657 (image[199],filter[1],mul_out[552][8]);
mul_8x8bit m1658 (image[200],filter[2],mul_out[552][9]);
mul_8x8bit m1659 (image[226],filter[3],mul_out[553][7]);
mul_8x8bit m1660 (image[227],filter[4],mul_out[553][8]);
mul_8x8bit m1661 (image[228],filter[5],mul_out[553][9]);
mul_8x8bit m1662 (image[254],filter[6],mul_out[554][7]);
mul_8x8bit m1663 (image[255],filter[7],mul_out[554][8]);
mul_8x8bit m1664 (image[256],filter[8],mul_out[554][9]);

adder_8bit ad184 (mul_out[552][7],mul_out[552][8],mul_out[552][9],mul_out[553][7],mul_out[553][8],mul_out[553][9],mul_out[554][7],mul_out[554][8],mul_out[554][9],conv_out[184]);



mul_8x8bit m1665 (image[199],filter[0],mul_out[555][7]);
mul_8x8bit m1666 (image[200],filter[1],mul_out[555][8]);
mul_8x8bit m1667 (image[201],filter[2],mul_out[555][9]);
mul_8x8bit m1668 (image[227],filter[3],mul_out[556][7]);
mul_8x8bit m1669 (image[228],filter[4],mul_out[556][8]);
mul_8x8bit m1670 (image[229],filter[5],mul_out[556][9]);
mul_8x8bit m1671 (image[255],filter[6],mul_out[557][7]);
mul_8x8bit m1672 (image[256],filter[7],mul_out[557][8]);
mul_8x8bit m1673 (image[257],filter[8],mul_out[557][9]);

adder_8bit ad185 (mul_out[555][7],mul_out[555][8],mul_out[555][9],mul_out[556][7],mul_out[556][8],mul_out[556][9],mul_out[557][7],mul_out[557][8],mul_out[557][9],conv_out[185]);



mul_8x8bit m1674 (image[200],filter[0],mul_out[558][7]);
mul_8x8bit m1675 (image[201],filter[1],mul_out[558][8]);
mul_8x8bit m1676 (image[202],filter[2],mul_out[558][9]);
mul_8x8bit m1677 (image[228],filter[3],mul_out[559][7]);
mul_8x8bit m1678 (image[229],filter[4],mul_out[559][8]);
mul_8x8bit m1679 (image[230],filter[5],mul_out[559][9]);
mul_8x8bit m1680 (image[256],filter[6],mul_out[560][7]);
mul_8x8bit m1681 (image[257],filter[7],mul_out[560][8]);
mul_8x8bit m1682 (image[258],filter[8],mul_out[560][9]);

adder_8bit ad186 (mul_out[558][7],mul_out[558][8],mul_out[558][9],mul_out[559][7],mul_out[559][8],mul_out[559][9],mul_out[560][7],mul_out[560][8],mul_out[560][9],conv_out[186]);



mul_8x8bit m1683 (image[201],filter[0],mul_out[561][7]);
mul_8x8bit m1684 (image[202],filter[1],mul_out[561][8]);
mul_8x8bit m1685 (image[203],filter[2],mul_out[561][9]);
mul_8x8bit m1686 (image[229],filter[3],mul_out[562][7]);
mul_8x8bit m1687 (image[230],filter[4],mul_out[562][8]);
mul_8x8bit m1688 (image[231],filter[5],mul_out[562][9]);
mul_8x8bit m1689 (image[257],filter[6],mul_out[563][7]);
mul_8x8bit m1690 (image[258],filter[7],mul_out[563][8]);
mul_8x8bit m1691 (image[259],filter[8],mul_out[563][9]);

adder_8bit ad187 (mul_out[561][7],mul_out[561][8],mul_out[561][9],mul_out[562][7],mul_out[562][8],mul_out[562][9],mul_out[563][7],mul_out[563][8],mul_out[563][9],conv_out[187]);



mul_8x8bit m1692 (image[202],filter[0],mul_out[564][7]);
mul_8x8bit m1693 (image[203],filter[1],mul_out[564][8]);
mul_8x8bit m1694 (image[204],filter[2],mul_out[564][9]);
mul_8x8bit m1695 (image[230],filter[3],mul_out[565][7]);
mul_8x8bit m1696 (image[231],filter[4],mul_out[565][8]);
mul_8x8bit m1697 (image[232],filter[5],mul_out[565][9]);
mul_8x8bit m1698 (image[258],filter[6],mul_out[566][7]);
mul_8x8bit m1699 (image[259],filter[7],mul_out[566][8]);
mul_8x8bit m1700 (image[260],filter[8],mul_out[566][9]);

adder_8bit ad188 (mul_out[564][7],mul_out[564][8],mul_out[564][9],mul_out[565][7],mul_out[565][8],mul_out[565][9],mul_out[566][7],mul_out[566][8],mul_out[566][9],conv_out[188]);



mul_8x8bit m1701 (image[203],filter[0],mul_out[567][7]);
mul_8x8bit m1702 (image[204],filter[1],mul_out[567][8]);
mul_8x8bit m1703 (image[205],filter[2],mul_out[567][9]);
mul_8x8bit m1704 (image[231],filter[3],mul_out[568][7]);
mul_8x8bit m1705 (image[232],filter[4],mul_out[568][8]);
mul_8x8bit m1706 (image[233],filter[5],mul_out[568][9]);
mul_8x8bit m1707 (image[259],filter[6],mul_out[569][7]);
mul_8x8bit m1708 (image[260],filter[7],mul_out[569][8]);
mul_8x8bit m1709 (image[261],filter[8],mul_out[569][9]);

adder_8bit ad189 (mul_out[567][7],mul_out[567][8],mul_out[567][9],mul_out[568][7],mul_out[568][8],mul_out[568][9],mul_out[569][7],mul_out[569][8],mul_out[569][9],conv_out[189]);



mul_8x8bit m1710 (image[204],filter[0],mul_out[570][7]);
mul_8x8bit m1711 (image[205],filter[1],mul_out[570][8]);
mul_8x8bit m1712 (image[206],filter[2],mul_out[570][9]);
mul_8x8bit m1713 (image[232],filter[3],mul_out[571][7]);
mul_8x8bit m1714 (image[233],filter[4],mul_out[571][8]);
mul_8x8bit m1715 (image[234],filter[5],mul_out[571][9]);
mul_8x8bit m1716 (image[260],filter[6],mul_out[572][7]);
mul_8x8bit m1717 (image[261],filter[7],mul_out[572][8]);
mul_8x8bit m1718 (image[262],filter[8],mul_out[572][9]);

adder_8bit ad190 (mul_out[570][7],mul_out[570][8],mul_out[570][9],mul_out[571][7],mul_out[571][8],mul_out[571][9],mul_out[572][7],mul_out[572][8],mul_out[572][9],conv_out[190]);



mul_8x8bit m1719 (image[205],filter[0],mul_out[573][7]);
mul_8x8bit m1720 (image[206],filter[1],mul_out[573][8]);
mul_8x8bit m1721 (image[207],filter[2],mul_out[573][9]);
mul_8x8bit m1722 (image[233],filter[3],mul_out[574][7]);
mul_8x8bit m1723 (image[234],filter[4],mul_out[574][8]);
mul_8x8bit m1724 (image[235],filter[5],mul_out[574][9]);
mul_8x8bit m1725 (image[261],filter[6],mul_out[575][7]);
mul_8x8bit m1726 (image[262],filter[7],mul_out[575][8]);
mul_8x8bit m1727 (image[263],filter[8],mul_out[575][9]);

adder_8bit ad191 (mul_out[573][7],mul_out[573][8],mul_out[573][9],mul_out[574][7],mul_out[574][8],mul_out[574][9],mul_out[575][7],mul_out[575][8],mul_out[575][9],conv_out[191]);



mul_8x8bit m1728 (image[206],filter[0],mul_out[576][7]);
mul_8x8bit m1729 (image[207],filter[1],mul_out[576][8]);
mul_8x8bit m1730 (image[208],filter[2],mul_out[576][9]);
mul_8x8bit m1731 (image[234],filter[3],mul_out[577][7]);
mul_8x8bit m1732 (image[235],filter[4],mul_out[577][8]);
mul_8x8bit m1733 (image[236],filter[5],mul_out[577][9]);
mul_8x8bit m1734 (image[262],filter[6],mul_out[578][7]);
mul_8x8bit m1735 (image[263],filter[7],mul_out[578][8]);
mul_8x8bit m1736 (image[264],filter[8],mul_out[578][9]);

adder_8bit ad192 (mul_out[576][7],mul_out[576][8],mul_out[576][9],mul_out[577][7],mul_out[577][8],mul_out[577][9],mul_out[578][7],mul_out[578][8],mul_out[578][9],conv_out[192]);



mul_8x8bit m1737 (image[207],filter[0],mul_out[579][7]);
mul_8x8bit m1738 (image[208],filter[1],mul_out[579][8]);
mul_8x8bit m1739 (image[209],filter[2],mul_out[579][9]);
mul_8x8bit m1740 (image[235],filter[3],mul_out[580][7]);
mul_8x8bit m1741 (image[236],filter[4],mul_out[580][8]);
mul_8x8bit m1742 (image[237],filter[5],mul_out[580][9]);
mul_8x8bit m1743 (image[263],filter[6],mul_out[581][7]);
mul_8x8bit m1744 (image[264],filter[7],mul_out[581][8]);
mul_8x8bit m1745 (image[265],filter[8],mul_out[581][9]);

adder_8bit ad193 (mul_out[579][7],mul_out[579][8],mul_out[579][9],mul_out[580][7],mul_out[580][8],mul_out[580][9],mul_out[581][7],mul_out[581][8],mul_out[581][9],conv_out[193]);



mul_8x8bit m1746 (image[208],filter[0],mul_out[582][7]);
mul_8x8bit m1747 (image[209],filter[1],mul_out[582][8]);
mul_8x8bit m1748 (image[210],filter[2],mul_out[582][9]);
mul_8x8bit m1749 (image[236],filter[3],mul_out[583][7]);
mul_8x8bit m1750 (image[237],filter[4],mul_out[583][8]);
mul_8x8bit m1751 (image[238],filter[5],mul_out[583][9]);
mul_8x8bit m1752 (image[264],filter[6],mul_out[584][7]);
mul_8x8bit m1753 (image[265],filter[7],mul_out[584][8]);
mul_8x8bit m1754 (image[266],filter[8],mul_out[584][9]);

adder_8bit ad194 (mul_out[582][7],mul_out[582][8],mul_out[582][9],mul_out[583][7],mul_out[583][8],mul_out[583][9],mul_out[584][7],mul_out[584][8],mul_out[584][9],conv_out[194]);



mul_8x8bit m1755 (image[209],filter[0],mul_out[585][7]);
mul_8x8bit m1756 (image[210],filter[1],mul_out[585][8]);
mul_8x8bit m1757 (image[211],filter[2],mul_out[585][9]);
mul_8x8bit m1758 (image[237],filter[3],mul_out[586][7]);
mul_8x8bit m1759 (image[238],filter[4],mul_out[586][8]);
mul_8x8bit m1760 (image[239],filter[5],mul_out[586][9]);
mul_8x8bit m1761 (image[265],filter[6],mul_out[587][7]);
mul_8x8bit m1762 (image[266],filter[7],mul_out[587][8]);
mul_8x8bit m1763 (image[267],filter[8],mul_out[587][9]);

adder_8bit ad195 (mul_out[585][7],mul_out[585][8],mul_out[585][9],mul_out[586][7],mul_out[586][8],mul_out[586][9],mul_out[587][7],mul_out[587][8],mul_out[587][9],conv_out[195]);



mul_8x8bit m1764 (image[210],filter[0],mul_out[588][7]);
mul_8x8bit m1765 (image[211],filter[1],mul_out[588][8]);
mul_8x8bit m1766 (image[212],filter[2],mul_out[588][9]);
mul_8x8bit m1767 (image[238],filter[3],mul_out[589][7]);
mul_8x8bit m1768 (image[239],filter[4],mul_out[589][8]);
mul_8x8bit m1769 (image[240],filter[5],mul_out[589][9]);
mul_8x8bit m1770 (image[266],filter[6],mul_out[590][7]);
mul_8x8bit m1771 (image[267],filter[7],mul_out[590][8]);
mul_8x8bit m1772 (image[268],filter[8],mul_out[590][9]);

adder_8bit ad196 (mul_out[588][7],mul_out[588][8],mul_out[588][9],mul_out[589][7],mul_out[589][8],mul_out[589][9],mul_out[590][7],mul_out[590][8],mul_out[590][9],conv_out[196]);



mul_8x8bit m1773 (image[211],filter[0],mul_out[591][7]);
mul_8x8bit m1774 (image[212],filter[1],mul_out[591][8]);
mul_8x8bit m1775 (image[213],filter[2],mul_out[591][9]);
mul_8x8bit m1776 (image[239],filter[3],mul_out[592][7]);
mul_8x8bit m1777 (image[240],filter[4],mul_out[592][8]);
mul_8x8bit m1778 (image[241],filter[5],mul_out[592][9]);
mul_8x8bit m1779 (image[267],filter[6],mul_out[593][7]);
mul_8x8bit m1780 (image[268],filter[7],mul_out[593][8]);
mul_8x8bit m1781 (image[269],filter[8],mul_out[593][9]);

adder_8bit ad197 (mul_out[591][7],mul_out[591][8],mul_out[591][9],mul_out[592][7],mul_out[592][8],mul_out[592][9],mul_out[593][7],mul_out[593][8],mul_out[593][9],conv_out[197]);



mul_8x8bit m1782 (image[212],filter[0],mul_out[594][7]);
mul_8x8bit m1783 (image[213],filter[1],mul_out[594][8]);
mul_8x8bit m1784 (image[214],filter[2],mul_out[594][9]);
mul_8x8bit m1785 (image[240],filter[3],mul_out[595][7]);
mul_8x8bit m1786 (image[241],filter[4],mul_out[595][8]);
mul_8x8bit m1787 (image[242],filter[5],mul_out[595][9]);
mul_8x8bit m1788 (image[268],filter[6],mul_out[596][7]);
mul_8x8bit m1789 (image[269],filter[7],mul_out[596][8]);
mul_8x8bit m1790 (image[270],filter[8],mul_out[596][9]);

adder_8bit ad198 (mul_out[594][7],mul_out[594][8],mul_out[594][9],mul_out[595][7],mul_out[595][8],mul_out[595][9],mul_out[596][7],mul_out[596][8],mul_out[596][9],conv_out[198]);



mul_8x8bit m1791 (image[213],filter[0],mul_out[597][7]);
mul_8x8bit m1792 (image[214],filter[1],mul_out[597][8]);
mul_8x8bit m1793 (image[215],filter[2],mul_out[597][9]);
mul_8x8bit m1794 (image[241],filter[3],mul_out[598][7]);
mul_8x8bit m1795 (image[242],filter[4],mul_out[598][8]);
mul_8x8bit m1796 (image[243],filter[5],mul_out[598][9]);
mul_8x8bit m1797 (image[269],filter[6],mul_out[599][7]);
mul_8x8bit m1798 (image[270],filter[7],mul_out[599][8]);
mul_8x8bit m1799 (image[271],filter[8],mul_out[599][9]);

adder_8bit ad199 (mul_out[597][7],mul_out[597][8],mul_out[597][9],mul_out[598][7],mul_out[598][8],mul_out[598][9],mul_out[599][7],mul_out[599][8],mul_out[599][9],conv_out[199]);



mul_8x8bit m1800 (image[214],filter[0],mul_out[600][7]);
mul_8x8bit m1801 (image[215],filter[1],mul_out[600][8]);
mul_8x8bit m1802 (image[216],filter[2],mul_out[600][9]);
mul_8x8bit m1803 (image[242],filter[3],mul_out[601][7]);
mul_8x8bit m1804 (image[243],filter[4],mul_out[601][8]);
mul_8x8bit m1805 (image[244],filter[5],mul_out[601][9]);
mul_8x8bit m1806 (image[270],filter[6],mul_out[602][7]);
mul_8x8bit m1807 (image[271],filter[7],mul_out[602][8]);
mul_8x8bit m1808 (image[272],filter[8],mul_out[602][9]);

adder_8bit ad200 (mul_out[600][7],mul_out[600][8],mul_out[600][9],mul_out[601][7],mul_out[601][8],mul_out[601][9],mul_out[602][7],mul_out[602][8],mul_out[602][9],conv_out[200]);



mul_8x8bit m1809 (image[215],filter[0],mul_out[603][7]);
mul_8x8bit m1810 (image[216],filter[1],mul_out[603][8]);
mul_8x8bit m1811 (image[217],filter[2],mul_out[603][9]);
mul_8x8bit m1812 (image[243],filter[3],mul_out[604][7]);
mul_8x8bit m1813 (image[244],filter[4],mul_out[604][8]);
mul_8x8bit m1814 (image[245],filter[5],mul_out[604][9]);
mul_8x8bit m1815 (image[271],filter[6],mul_out[605][7]);
mul_8x8bit m1816 (image[272],filter[7],mul_out[605][8]);
mul_8x8bit m1817 (image[273],filter[8],mul_out[605][9]);

adder_8bit ad201 (mul_out[603][7],mul_out[603][8],mul_out[603][9],mul_out[604][7],mul_out[604][8],mul_out[604][9],mul_out[605][7],mul_out[605][8],mul_out[605][9],conv_out[201]);



mul_8x8bit m1818 (image[216],filter[0],mul_out[606][7]);
mul_8x8bit m1819 (image[217],filter[1],mul_out[606][8]);
mul_8x8bit m1820 (image[218],filter[2],mul_out[606][9]);
mul_8x8bit m1821 (image[244],filter[3],mul_out[607][7]);
mul_8x8bit m1822 (image[245],filter[4],mul_out[607][8]);
mul_8x8bit m1823 (image[246],filter[5],mul_out[607][9]);
mul_8x8bit m1824 (image[272],filter[6],mul_out[608][7]);
mul_8x8bit m1825 (image[273],filter[7],mul_out[608][8]);
mul_8x8bit m1826 (image[274],filter[8],mul_out[608][9]);

adder_8bit ad202 (mul_out[606][7],mul_out[606][8],mul_out[606][9],mul_out[607][7],mul_out[607][8],mul_out[607][9],mul_out[608][7],mul_out[608][8],mul_out[608][9],conv_out[202]);



mul_8x8bit m1827 (image[217],filter[0],mul_out[609][7]);
mul_8x8bit m1828 (image[218],filter[1],mul_out[609][8]);
mul_8x8bit m1829 (image[219],filter[2],mul_out[609][9]);
mul_8x8bit m1830 (image[245],filter[3],mul_out[610][7]);
mul_8x8bit m1831 (image[246],filter[4],mul_out[610][8]);
mul_8x8bit m1832 (image[247],filter[5],mul_out[610][9]);
mul_8x8bit m1833 (image[273],filter[6],mul_out[611][7]);
mul_8x8bit m1834 (image[274],filter[7],mul_out[611][8]);
mul_8x8bit m1835 (image[275],filter[8],mul_out[611][9]);

adder_8bit ad203 (mul_out[609][7],mul_out[609][8],mul_out[609][9],mul_out[610][7],mul_out[610][8],mul_out[610][9],mul_out[611][7],mul_out[611][8],mul_out[611][9],conv_out[203]);



mul_8x8bit m1836 (image[218],filter[0],mul_out[612][7]);
mul_8x8bit m1837 (image[219],filter[1],mul_out[612][8]);
mul_8x8bit m1838 (image[220],filter[2],mul_out[612][9]);
mul_8x8bit m1839 (image[246],filter[3],mul_out[613][7]);
mul_8x8bit m1840 (image[247],filter[4],mul_out[613][8]);
mul_8x8bit m1841 (image[248],filter[5],mul_out[613][9]);
mul_8x8bit m1842 (image[274],filter[6],mul_out[614][7]);
mul_8x8bit m1843 (image[275],filter[7],mul_out[614][8]);
mul_8x8bit m1844 (image[276],filter[8],mul_out[614][9]);

adder_8bit ad204 (mul_out[612][7],mul_out[612][8],mul_out[612][9],mul_out[613][7],mul_out[613][8],mul_out[613][9],mul_out[614][7],mul_out[614][8],mul_out[614][9],conv_out[204]);



mul_8x8bit m1845 (image[219],filter[0],mul_out[615][7]);
mul_8x8bit m1846 (image[220],filter[1],mul_out[615][8]);
mul_8x8bit m1847 (image[221],filter[2],mul_out[615][9]);
mul_8x8bit m1848 (image[247],filter[3],mul_out[616][7]);
mul_8x8bit m1849 (image[248],filter[4],mul_out[616][8]);
mul_8x8bit m1850 (image[249],filter[5],mul_out[616][9]);
mul_8x8bit m1851 (image[275],filter[6],mul_out[617][7]);
mul_8x8bit m1852 (image[276],filter[7],mul_out[617][8]);
mul_8x8bit m1853 (image[277],filter[8],mul_out[617][9]);

adder_8bit ad205 (mul_out[615][7],mul_out[615][8],mul_out[615][9],mul_out[616][7],mul_out[616][8],mul_out[616][9],mul_out[617][7],mul_out[617][8],mul_out[617][9],conv_out[205]);



mul_8x8bit m1854 (image[220],filter[0],mul_out[618][7]);
mul_8x8bit m1855 (image[221],filter[1],mul_out[618][8]);
mul_8x8bit m1856 (image[222],filter[2],mul_out[618][9]);
mul_8x8bit m1857 (image[248],filter[3],mul_out[619][7]);
mul_8x8bit m1858 (image[249],filter[4],mul_out[619][8]);
mul_8x8bit m1859 (image[250],filter[5],mul_out[619][9]);
mul_8x8bit m1860 (image[276],filter[6],mul_out[620][7]);
mul_8x8bit m1861 (image[277],filter[7],mul_out[620][8]);
mul_8x8bit m1862 (image[278],filter[8],mul_out[620][9]);

adder_8bit ad206 (mul_out[618][7],mul_out[618][8],mul_out[618][9],mul_out[619][7],mul_out[619][8],mul_out[619][9],mul_out[620][7],mul_out[620][8],mul_out[620][9],conv_out[206]);



mul_8x8bit m1863 (image[221],filter[0],mul_out[621][7]);
mul_8x8bit m1864 (image[222],filter[1],mul_out[621][8]);
mul_8x8bit m1865 (image[223],filter[2],mul_out[621][9]);
mul_8x8bit m1866 (image[249],filter[3],mul_out[622][7]);
mul_8x8bit m1867 (image[250],filter[4],mul_out[622][8]);
mul_8x8bit m1868 (image[251],filter[5],mul_out[622][9]);
mul_8x8bit m1869 (image[277],filter[6],mul_out[623][7]);
mul_8x8bit m1870 (image[278],filter[7],mul_out[623][8]);
mul_8x8bit m1871 (image[279],filter[8],mul_out[623][9]);

adder_8bit ad207 (mul_out[621][7],mul_out[621][8],mul_out[621][9],mul_out[622][7],mul_out[622][8],mul_out[622][9],mul_out[623][7],mul_out[623][8],mul_out[623][9],conv_out[207]);



mul_8x8bit m1872 (image[224],filter[0],mul_out[624][8]);
mul_8x8bit m1873 (image[225],filter[1],mul_out[624][9]);
mul_8x8bit m1874 (image[226],filter[2],mul_out[624][10]);
mul_8x8bit m1875 (image[252],filter[3],mul_out[625][8]);
mul_8x8bit m1876 (image[253],filter[4],mul_out[625][9]);
mul_8x8bit m1877 (image[254],filter[5],mul_out[625][10]);
mul_8x8bit m1878 (image[280],filter[6],mul_out[626][8]);
mul_8x8bit m1879 (image[281],filter[7],mul_out[626][9]);
mul_8x8bit m1880 (image[282],filter[8],mul_out[626][10]);

adder_8bit ad208 (mul_out[624][8],mul_out[624][9],mul_out[624][10],mul_out[625][8],mul_out[625][9],mul_out[625][10],mul_out[626][8],mul_out[626][9],mul_out[626][10],conv_out[208]);



mul_8x8bit m1881 (image[225],filter[0],mul_out[627][8]);
mul_8x8bit m1882 (image[226],filter[1],mul_out[627][9]);
mul_8x8bit m1883 (image[227],filter[2],mul_out[627][10]);
mul_8x8bit m1884 (image[253],filter[3],mul_out[628][8]);
mul_8x8bit m1885 (image[254],filter[4],mul_out[628][9]);
mul_8x8bit m1886 (image[255],filter[5],mul_out[628][10]);
mul_8x8bit m1887 (image[281],filter[6],mul_out[629][8]);
mul_8x8bit m1888 (image[282],filter[7],mul_out[629][9]);
mul_8x8bit m1889 (image[283],filter[8],mul_out[629][10]);

adder_8bit ad209 (mul_out[627][8],mul_out[627][9],mul_out[627][10],mul_out[628][8],mul_out[628][9],mul_out[628][10],mul_out[629][8],mul_out[629][9],mul_out[629][10],conv_out[209]);



mul_8x8bit m1890 (image[226],filter[0],mul_out[630][8]);
mul_8x8bit m1891 (image[227],filter[1],mul_out[630][9]);
mul_8x8bit m1892 (image[228],filter[2],mul_out[630][10]);
mul_8x8bit m1893 (image[254],filter[3],mul_out[631][8]);
mul_8x8bit m1894 (image[255],filter[4],mul_out[631][9]);
mul_8x8bit m1895 (image[256],filter[5],mul_out[631][10]);
mul_8x8bit m1896 (image[282],filter[6],mul_out[632][8]);
mul_8x8bit m1897 (image[283],filter[7],mul_out[632][9]);
mul_8x8bit m1898 (image[284],filter[8],mul_out[632][10]);

adder_8bit ad210 (mul_out[630][8],mul_out[630][9],mul_out[630][10],mul_out[631][8],mul_out[631][9],mul_out[631][10],mul_out[632][8],mul_out[632][9],mul_out[632][10],conv_out[210]);



mul_8x8bit m1899 (image[227],filter[0],mul_out[633][8]);
mul_8x8bit m1900 (image[228],filter[1],mul_out[633][9]);
mul_8x8bit m1901 (image[229],filter[2],mul_out[633][10]);
mul_8x8bit m1902 (image[255],filter[3],mul_out[634][8]);
mul_8x8bit m1903 (image[256],filter[4],mul_out[634][9]);
mul_8x8bit m1904 (image[257],filter[5],mul_out[634][10]);
mul_8x8bit m1905 (image[283],filter[6],mul_out[635][8]);
mul_8x8bit m1906 (image[284],filter[7],mul_out[635][9]);
mul_8x8bit m1907 (image[285],filter[8],mul_out[635][10]);

adder_8bit ad211 (mul_out[633][8],mul_out[633][9],mul_out[633][10],mul_out[634][8],mul_out[634][9],mul_out[634][10],mul_out[635][8],mul_out[635][9],mul_out[635][10],conv_out[211]);



mul_8x8bit m1908 (image[228],filter[0],mul_out[636][8]);
mul_8x8bit m1909 (image[229],filter[1],mul_out[636][9]);
mul_8x8bit m1910 (image[230],filter[2],mul_out[636][10]);
mul_8x8bit m1911 (image[256],filter[3],mul_out[637][8]);
mul_8x8bit m1912 (image[257],filter[4],mul_out[637][9]);
mul_8x8bit m1913 (image[258],filter[5],mul_out[637][10]);
mul_8x8bit m1914 (image[284],filter[6],mul_out[638][8]);
mul_8x8bit m1915 (image[285],filter[7],mul_out[638][9]);
mul_8x8bit m1916 (image[286],filter[8],mul_out[638][10]);

adder_8bit ad212 (mul_out[636][8],mul_out[636][9],mul_out[636][10],mul_out[637][8],mul_out[637][9],mul_out[637][10],mul_out[638][8],mul_out[638][9],mul_out[638][10],conv_out[212]);



mul_8x8bit m1917 (image[229],filter[0],mul_out[639][8]);
mul_8x8bit m1918 (image[230],filter[1],mul_out[639][9]);
mul_8x8bit m1919 (image[231],filter[2],mul_out[639][10]);
mul_8x8bit m1920 (image[257],filter[3],mul_out[640][8]);
mul_8x8bit m1921 (image[258],filter[4],mul_out[640][9]);
mul_8x8bit m1922 (image[259],filter[5],mul_out[640][10]);
mul_8x8bit m1923 (image[285],filter[6],mul_out[641][8]);
mul_8x8bit m1924 (image[286],filter[7],mul_out[641][9]);
mul_8x8bit m1925 (image[287],filter[8],mul_out[641][10]);

adder_8bit ad213 (mul_out[639][8],mul_out[639][9],mul_out[639][10],mul_out[640][8],mul_out[640][9],mul_out[640][10],mul_out[641][8],mul_out[641][9],mul_out[641][10],conv_out[213]);



mul_8x8bit m1926 (image[230],filter[0],mul_out[642][8]);
mul_8x8bit m1927 (image[231],filter[1],mul_out[642][9]);
mul_8x8bit m1928 (image[232],filter[2],mul_out[642][10]);
mul_8x8bit m1929 (image[258],filter[3],mul_out[643][8]);
mul_8x8bit m1930 (image[259],filter[4],mul_out[643][9]);
mul_8x8bit m1931 (image[260],filter[5],mul_out[643][10]);
mul_8x8bit m1932 (image[286],filter[6],mul_out[644][8]);
mul_8x8bit m1933 (image[287],filter[7],mul_out[644][9]);
mul_8x8bit m1934 (image[288],filter[8],mul_out[644][10]);

adder_8bit ad214 (mul_out[642][8],mul_out[642][9],mul_out[642][10],mul_out[643][8],mul_out[643][9],mul_out[643][10],mul_out[644][8],mul_out[644][9],mul_out[644][10],conv_out[214]);



mul_8x8bit m1935 (image[231],filter[0],mul_out[645][8]);
mul_8x8bit m1936 (image[232],filter[1],mul_out[645][9]);
mul_8x8bit m1937 (image[233],filter[2],mul_out[645][10]);
mul_8x8bit m1938 (image[259],filter[3],mul_out[646][8]);
mul_8x8bit m1939 (image[260],filter[4],mul_out[646][9]);
mul_8x8bit m1940 (image[261],filter[5],mul_out[646][10]);
mul_8x8bit m1941 (image[287],filter[6],mul_out[647][8]);
mul_8x8bit m1942 (image[288],filter[7],mul_out[647][9]);
mul_8x8bit m1943 (image[289],filter[8],mul_out[647][10]);

adder_8bit ad215 (mul_out[645][8],mul_out[645][9],mul_out[645][10],mul_out[646][8],mul_out[646][9],mul_out[646][10],mul_out[647][8],mul_out[647][9],mul_out[647][10],conv_out[215]);



mul_8x8bit m1944 (image[232],filter[0],mul_out[648][8]);
mul_8x8bit m1945 (image[233],filter[1],mul_out[648][9]);
mul_8x8bit m1946 (image[234],filter[2],mul_out[648][10]);
mul_8x8bit m1947 (image[260],filter[3],mul_out[649][8]);
mul_8x8bit m1948 (image[261],filter[4],mul_out[649][9]);
mul_8x8bit m1949 (image[262],filter[5],mul_out[649][10]);
mul_8x8bit m1950 (image[288],filter[6],mul_out[650][8]);
mul_8x8bit m1951 (image[289],filter[7],mul_out[650][9]);
mul_8x8bit m1952 (image[290],filter[8],mul_out[650][10]);

adder_8bit ad216 (mul_out[648][8],mul_out[648][9],mul_out[648][10],mul_out[649][8],mul_out[649][9],mul_out[649][10],mul_out[650][8],mul_out[650][9],mul_out[650][10],conv_out[216]);



mul_8x8bit m1953 (image[233],filter[0],mul_out[651][8]);
mul_8x8bit m1954 (image[234],filter[1],mul_out[651][9]);
mul_8x8bit m1955 (image[235],filter[2],mul_out[651][10]);
mul_8x8bit m1956 (image[261],filter[3],mul_out[652][8]);
mul_8x8bit m1957 (image[262],filter[4],mul_out[652][9]);
mul_8x8bit m1958 (image[263],filter[5],mul_out[652][10]);
mul_8x8bit m1959 (image[289],filter[6],mul_out[653][8]);
mul_8x8bit m1960 (image[290],filter[7],mul_out[653][9]);
mul_8x8bit m1961 (image[291],filter[8],mul_out[653][10]);

adder_8bit ad217 (mul_out[651][8],mul_out[651][9],mul_out[651][10],mul_out[652][8],mul_out[652][9],mul_out[652][10],mul_out[653][8],mul_out[653][9],mul_out[653][10],conv_out[217]);



mul_8x8bit m1962 (image[234],filter[0],mul_out[654][8]);
mul_8x8bit m1963 (image[235],filter[1],mul_out[654][9]);
mul_8x8bit m1964 (image[236],filter[2],mul_out[654][10]);
mul_8x8bit m1965 (image[262],filter[3],mul_out[655][8]);
mul_8x8bit m1966 (image[263],filter[4],mul_out[655][9]);
mul_8x8bit m1967 (image[264],filter[5],mul_out[655][10]);
mul_8x8bit m1968 (image[290],filter[6],mul_out[656][8]);
mul_8x8bit m1969 (image[291],filter[7],mul_out[656][9]);
mul_8x8bit m1970 (image[292],filter[8],mul_out[656][10]);

adder_8bit ad218 (mul_out[654][8],mul_out[654][9],mul_out[654][10],mul_out[655][8],mul_out[655][9],mul_out[655][10],mul_out[656][8],mul_out[656][9],mul_out[656][10],conv_out[218]);



mul_8x8bit m1971 (image[235],filter[0],mul_out[657][8]);
mul_8x8bit m1972 (image[236],filter[1],mul_out[657][9]);
mul_8x8bit m1973 (image[237],filter[2],mul_out[657][10]);
mul_8x8bit m1974 (image[263],filter[3],mul_out[658][8]);
mul_8x8bit m1975 (image[264],filter[4],mul_out[658][9]);
mul_8x8bit m1976 (image[265],filter[5],mul_out[658][10]);
mul_8x8bit m1977 (image[291],filter[6],mul_out[659][8]);
mul_8x8bit m1978 (image[292],filter[7],mul_out[659][9]);
mul_8x8bit m1979 (image[293],filter[8],mul_out[659][10]);

adder_8bit ad219 (mul_out[657][8],mul_out[657][9],mul_out[657][10],mul_out[658][8],mul_out[658][9],mul_out[658][10],mul_out[659][8],mul_out[659][9],mul_out[659][10],conv_out[219]);



mul_8x8bit m1980 (image[236],filter[0],mul_out[660][8]);
mul_8x8bit m1981 (image[237],filter[1],mul_out[660][9]);
mul_8x8bit m1982 (image[238],filter[2],mul_out[660][10]);
mul_8x8bit m1983 (image[264],filter[3],mul_out[661][8]);
mul_8x8bit m1984 (image[265],filter[4],mul_out[661][9]);
mul_8x8bit m1985 (image[266],filter[5],mul_out[661][10]);
mul_8x8bit m1986 (image[292],filter[6],mul_out[662][8]);
mul_8x8bit m1987 (image[293],filter[7],mul_out[662][9]);
mul_8x8bit m1988 (image[294],filter[8],mul_out[662][10]);

adder_8bit ad220 (mul_out[660][8],mul_out[660][9],mul_out[660][10],mul_out[661][8],mul_out[661][9],mul_out[661][10],mul_out[662][8],mul_out[662][9],mul_out[662][10],conv_out[220]);



mul_8x8bit m1989 (image[237],filter[0],mul_out[663][8]);
mul_8x8bit m1990 (image[238],filter[1],mul_out[663][9]);
mul_8x8bit m1991 (image[239],filter[2],mul_out[663][10]);
mul_8x8bit m1992 (image[265],filter[3],mul_out[664][8]);
mul_8x8bit m1993 (image[266],filter[4],mul_out[664][9]);
mul_8x8bit m1994 (image[267],filter[5],mul_out[664][10]);
mul_8x8bit m1995 (image[293],filter[6],mul_out[665][8]);
mul_8x8bit m1996 (image[294],filter[7],mul_out[665][9]);
mul_8x8bit m1997 (image[295],filter[8],mul_out[665][10]);

adder_8bit ad221 (mul_out[663][8],mul_out[663][9],mul_out[663][10],mul_out[664][8],mul_out[664][9],mul_out[664][10],mul_out[665][8],mul_out[665][9],mul_out[665][10],conv_out[221]);



mul_8x8bit m1998 (image[238],filter[0],mul_out[666][8]);
mul_8x8bit m1999 (image[239],filter[1],mul_out[666][9]);
mul_8x8bit m2000 (image[240],filter[2],mul_out[666][10]);
mul_8x8bit m2001 (image[266],filter[3],mul_out[667][8]);
mul_8x8bit m2002 (image[267],filter[4],mul_out[667][9]);
mul_8x8bit m2003 (image[268],filter[5],mul_out[667][10]);
mul_8x8bit m2004 (image[294],filter[6],mul_out[668][8]);
mul_8x8bit m2005 (image[295],filter[7],mul_out[668][9]);
mul_8x8bit m2006 (image[296],filter[8],mul_out[668][10]);

adder_8bit ad222 (mul_out[666][8],mul_out[666][9],mul_out[666][10],mul_out[667][8],mul_out[667][9],mul_out[667][10],mul_out[668][8],mul_out[668][9],mul_out[668][10],conv_out[222]);



mul_8x8bit m2007 (image[239],filter[0],mul_out[669][8]);
mul_8x8bit m2008 (image[240],filter[1],mul_out[669][9]);
mul_8x8bit m2009 (image[241],filter[2],mul_out[669][10]);
mul_8x8bit m2010 (image[267],filter[3],mul_out[670][8]);
mul_8x8bit m2011 (image[268],filter[4],mul_out[670][9]);
mul_8x8bit m2012 (image[269],filter[5],mul_out[670][10]);
mul_8x8bit m2013 (image[295],filter[6],mul_out[671][8]);
mul_8x8bit m2014 (image[296],filter[7],mul_out[671][9]);
mul_8x8bit m2015 (image[297],filter[8],mul_out[671][10]);

adder_8bit ad223 (mul_out[669][8],mul_out[669][9],mul_out[669][10],mul_out[670][8],mul_out[670][9],mul_out[670][10],mul_out[671][8],mul_out[671][9],mul_out[671][10],conv_out[223]);



mul_8x8bit m2016 (image[240],filter[0],mul_out[672][8]);
mul_8x8bit m2017 (image[241],filter[1],mul_out[672][9]);
mul_8x8bit m2018 (image[242],filter[2],mul_out[672][10]);
mul_8x8bit m2019 (image[268],filter[3],mul_out[673][8]);
mul_8x8bit m2020 (image[269],filter[4],mul_out[673][9]);
mul_8x8bit m2021 (image[270],filter[5],mul_out[673][10]);
mul_8x8bit m2022 (image[296],filter[6],mul_out[674][8]);
mul_8x8bit m2023 (image[297],filter[7],mul_out[674][9]);
mul_8x8bit m2024 (image[298],filter[8],mul_out[674][10]);

adder_8bit ad224 (mul_out[672][8],mul_out[672][9],mul_out[672][10],mul_out[673][8],mul_out[673][9],mul_out[673][10],mul_out[674][8],mul_out[674][9],mul_out[674][10],conv_out[224]);



mul_8x8bit m2025 (image[241],filter[0],mul_out[675][8]);
mul_8x8bit m2026 (image[242],filter[1],mul_out[675][9]);
mul_8x8bit m2027 (image[243],filter[2],mul_out[675][10]);
mul_8x8bit m2028 (image[269],filter[3],mul_out[676][8]);
mul_8x8bit m2029 (image[270],filter[4],mul_out[676][9]);
mul_8x8bit m2030 (image[271],filter[5],mul_out[676][10]);
mul_8x8bit m2031 (image[297],filter[6],mul_out[677][8]);
mul_8x8bit m2032 (image[298],filter[7],mul_out[677][9]);
mul_8x8bit m2033 (image[299],filter[8],mul_out[677][10]);

adder_8bit ad225 (mul_out[675][8],mul_out[675][9],mul_out[675][10],mul_out[676][8],mul_out[676][9],mul_out[676][10],mul_out[677][8],mul_out[677][9],mul_out[677][10],conv_out[225]);



mul_8x8bit m2034 (image[242],filter[0],mul_out[678][8]);
mul_8x8bit m2035 (image[243],filter[1],mul_out[678][9]);
mul_8x8bit m2036 (image[244],filter[2],mul_out[678][10]);
mul_8x8bit m2037 (image[270],filter[3],mul_out[679][8]);
mul_8x8bit m2038 (image[271],filter[4],mul_out[679][9]);
mul_8x8bit m2039 (image[272],filter[5],mul_out[679][10]);
mul_8x8bit m2040 (image[298],filter[6],mul_out[680][8]);
mul_8x8bit m2041 (image[299],filter[7],mul_out[680][9]);
mul_8x8bit m2042 (image[300],filter[8],mul_out[680][10]);

adder_8bit ad226 (mul_out[678][8],mul_out[678][9],mul_out[678][10],mul_out[679][8],mul_out[679][9],mul_out[679][10],mul_out[680][8],mul_out[680][9],mul_out[680][10],conv_out[226]);



mul_8x8bit m2043 (image[243],filter[0],mul_out[681][8]);
mul_8x8bit m2044 (image[244],filter[1],mul_out[681][9]);
mul_8x8bit m2045 (image[245],filter[2],mul_out[681][10]);
mul_8x8bit m2046 (image[271],filter[3],mul_out[682][8]);
mul_8x8bit m2047 (image[272],filter[4],mul_out[682][9]);
mul_8x8bit m2048 (image[273],filter[5],mul_out[682][10]);
mul_8x8bit m2049 (image[299],filter[6],mul_out[683][8]);
mul_8x8bit m2050 (image[300],filter[7],mul_out[683][9]);
mul_8x8bit m2051 (image[301],filter[8],mul_out[683][10]);

adder_8bit ad227 (mul_out[681][8],mul_out[681][9],mul_out[681][10],mul_out[682][8],mul_out[682][9],mul_out[682][10],mul_out[683][8],mul_out[683][9],mul_out[683][10],conv_out[227]);



mul_8x8bit m2052 (image[244],filter[0],mul_out[684][8]);
mul_8x8bit m2053 (image[245],filter[1],mul_out[684][9]);
mul_8x8bit m2054 (image[246],filter[2],mul_out[684][10]);
mul_8x8bit m2055 (image[272],filter[3],mul_out[685][8]);
mul_8x8bit m2056 (image[273],filter[4],mul_out[685][9]);
mul_8x8bit m2057 (image[274],filter[5],mul_out[685][10]);
mul_8x8bit m2058 (image[300],filter[6],mul_out[686][8]);
mul_8x8bit m2059 (image[301],filter[7],mul_out[686][9]);
mul_8x8bit m2060 (image[302],filter[8],mul_out[686][10]);

adder_8bit ad228 (mul_out[684][8],mul_out[684][9],mul_out[684][10],mul_out[685][8],mul_out[685][9],mul_out[685][10],mul_out[686][8],mul_out[686][9],mul_out[686][10],conv_out[228]);



mul_8x8bit m2061 (image[245],filter[0],mul_out[687][8]);
mul_8x8bit m2062 (image[246],filter[1],mul_out[687][9]);
mul_8x8bit m2063 (image[247],filter[2],mul_out[687][10]);
mul_8x8bit m2064 (image[273],filter[3],mul_out[688][8]);
mul_8x8bit m2065 (image[274],filter[4],mul_out[688][9]);
mul_8x8bit m2066 (image[275],filter[5],mul_out[688][10]);
mul_8x8bit m2067 (image[301],filter[6],mul_out[689][8]);
mul_8x8bit m2068 (image[302],filter[7],mul_out[689][9]);
mul_8x8bit m2069 (image[303],filter[8],mul_out[689][10]);

adder_8bit ad229 (mul_out[687][8],mul_out[687][9],mul_out[687][10],mul_out[688][8],mul_out[688][9],mul_out[688][10],mul_out[689][8],mul_out[689][9],mul_out[689][10],conv_out[229]);



mul_8x8bit m2070 (image[246],filter[0],mul_out[690][8]);
mul_8x8bit m2071 (image[247],filter[1],mul_out[690][9]);
mul_8x8bit m2072 (image[248],filter[2],mul_out[690][10]);
mul_8x8bit m2073 (image[274],filter[3],mul_out[691][8]);
mul_8x8bit m2074 (image[275],filter[4],mul_out[691][9]);
mul_8x8bit m2075 (image[276],filter[5],mul_out[691][10]);
mul_8x8bit m2076 (image[302],filter[6],mul_out[692][8]);
mul_8x8bit m2077 (image[303],filter[7],mul_out[692][9]);
mul_8x8bit m2078 (image[304],filter[8],mul_out[692][10]);

adder_8bit ad230 (mul_out[690][8],mul_out[690][9],mul_out[690][10],mul_out[691][8],mul_out[691][9],mul_out[691][10],mul_out[692][8],mul_out[692][9],mul_out[692][10],conv_out[230]);



mul_8x8bit m2079 (image[247],filter[0],mul_out[693][8]);
mul_8x8bit m2080 (image[248],filter[1],mul_out[693][9]);
mul_8x8bit m2081 (image[249],filter[2],mul_out[693][10]);
mul_8x8bit m2082 (image[275],filter[3],mul_out[694][8]);
mul_8x8bit m2083 (image[276],filter[4],mul_out[694][9]);
mul_8x8bit m2084 (image[277],filter[5],mul_out[694][10]);
mul_8x8bit m2085 (image[303],filter[6],mul_out[695][8]);
mul_8x8bit m2086 (image[304],filter[7],mul_out[695][9]);
mul_8x8bit m2087 (image[305],filter[8],mul_out[695][10]);

adder_8bit ad231 (mul_out[693][8],mul_out[693][9],mul_out[693][10],mul_out[694][8],mul_out[694][9],mul_out[694][10],mul_out[695][8],mul_out[695][9],mul_out[695][10],conv_out[231]);



mul_8x8bit m2088 (image[248],filter[0],mul_out[696][8]);
mul_8x8bit m2089 (image[249],filter[1],mul_out[696][9]);
mul_8x8bit m2090 (image[250],filter[2],mul_out[696][10]);
mul_8x8bit m2091 (image[276],filter[3],mul_out[697][8]);
mul_8x8bit m2092 (image[277],filter[4],mul_out[697][9]);
mul_8x8bit m2093 (image[278],filter[5],mul_out[697][10]);
mul_8x8bit m2094 (image[304],filter[6],mul_out[698][8]);
mul_8x8bit m2095 (image[305],filter[7],mul_out[698][9]);
mul_8x8bit m2096 (image[306],filter[8],mul_out[698][10]);

adder_8bit ad232 (mul_out[696][8],mul_out[696][9],mul_out[696][10],mul_out[697][8],mul_out[697][9],mul_out[697][10],mul_out[698][8],mul_out[698][9],mul_out[698][10],conv_out[232]);



mul_8x8bit m2097 (image[249],filter[0],mul_out[699][8]);
mul_8x8bit m2098 (image[250],filter[1],mul_out[699][9]);
mul_8x8bit m2099 (image[251],filter[2],mul_out[699][10]);
mul_8x8bit m2100 (image[277],filter[3],mul_out[700][8]);
mul_8x8bit m2101 (image[278],filter[4],mul_out[700][9]);
mul_8x8bit m2102 (image[279],filter[5],mul_out[700][10]);
mul_8x8bit m2103 (image[305],filter[6],mul_out[701][8]);
mul_8x8bit m2104 (image[306],filter[7],mul_out[701][9]);
mul_8x8bit m2105 (image[307],filter[8],mul_out[701][10]);

adder_8bit ad233 (mul_out[699][8],mul_out[699][9],mul_out[699][10],mul_out[700][8],mul_out[700][9],mul_out[700][10],mul_out[701][8],mul_out[701][9],mul_out[701][10],conv_out[233]);



mul_8x8bit m2106 (image[252],filter[0],mul_out[702][9]);
mul_8x8bit m2107 (image[253],filter[1],mul_out[702][10]);
mul_8x8bit m2108 (image[254],filter[2],mul_out[702][11]);
mul_8x8bit m2109 (image[280],filter[3],mul_out[703][9]);
mul_8x8bit m2110 (image[281],filter[4],mul_out[703][10]);
mul_8x8bit m2111 (image[282],filter[5],mul_out[703][11]);
mul_8x8bit m2112 (image[308],filter[6],mul_out[704][9]);
mul_8x8bit m2113 (image[309],filter[7],mul_out[704][10]);
mul_8x8bit m2114 (image[310],filter[8],mul_out[704][11]);

adder_8bit ad234 (mul_out[702][9],mul_out[702][10],mul_out[702][11],mul_out[703][9],mul_out[703][10],mul_out[703][11],mul_out[704][9],mul_out[704][10],mul_out[704][11],conv_out[234]);



mul_8x8bit m2115 (image[253],filter[0],mul_out[705][9]);
mul_8x8bit m2116 (image[254],filter[1],mul_out[705][10]);
mul_8x8bit m2117 (image[255],filter[2],mul_out[705][11]);
mul_8x8bit m2118 (image[281],filter[3],mul_out[706][9]);
mul_8x8bit m2119 (image[282],filter[4],mul_out[706][10]);
mul_8x8bit m2120 (image[283],filter[5],mul_out[706][11]);
mul_8x8bit m2121 (image[309],filter[6],mul_out[707][9]);
mul_8x8bit m2122 (image[310],filter[7],mul_out[707][10]);
mul_8x8bit m2123 (image[311],filter[8],mul_out[707][11]);

adder_8bit ad235 (mul_out[705][9],mul_out[705][10],mul_out[705][11],mul_out[706][9],mul_out[706][10],mul_out[706][11],mul_out[707][9],mul_out[707][10],mul_out[707][11],conv_out[235]);



mul_8x8bit m2124 (image[254],filter[0],mul_out[708][9]);
mul_8x8bit m2125 (image[255],filter[1],mul_out[708][10]);
mul_8x8bit m2126 (image[256],filter[2],mul_out[708][11]);
mul_8x8bit m2127 (image[282],filter[3],mul_out[709][9]);
mul_8x8bit m2128 (image[283],filter[4],mul_out[709][10]);
mul_8x8bit m2129 (image[284],filter[5],mul_out[709][11]);
mul_8x8bit m2130 (image[310],filter[6],mul_out[710][9]);
mul_8x8bit m2131 (image[311],filter[7],mul_out[710][10]);
mul_8x8bit m2132 (image[312],filter[8],mul_out[710][11]);

adder_8bit ad236 (mul_out[708][9],mul_out[708][10],mul_out[708][11],mul_out[709][9],mul_out[709][10],mul_out[709][11],mul_out[710][9],mul_out[710][10],mul_out[710][11],conv_out[236]);



mul_8x8bit m2133 (image[255],filter[0],mul_out[711][9]);
mul_8x8bit m2134 (image[256],filter[1],mul_out[711][10]);
mul_8x8bit m2135 (image[257],filter[2],mul_out[711][11]);
mul_8x8bit m2136 (image[283],filter[3],mul_out[712][9]);
mul_8x8bit m2137 (image[284],filter[4],mul_out[712][10]);
mul_8x8bit m2138 (image[285],filter[5],mul_out[712][11]);
mul_8x8bit m2139 (image[311],filter[6],mul_out[713][9]);
mul_8x8bit m2140 (image[312],filter[7],mul_out[713][10]);
mul_8x8bit m2141 (image[313],filter[8],mul_out[713][11]);

adder_8bit ad237 (mul_out[711][9],mul_out[711][10],mul_out[711][11],mul_out[712][9],mul_out[712][10],mul_out[712][11],mul_out[713][9],mul_out[713][10],mul_out[713][11],conv_out[237]);



mul_8x8bit m2142 (image[256],filter[0],mul_out[714][9]);
mul_8x8bit m2143 (image[257],filter[1],mul_out[714][10]);
mul_8x8bit m2144 (image[258],filter[2],mul_out[714][11]);
mul_8x8bit m2145 (image[284],filter[3],mul_out[715][9]);
mul_8x8bit m2146 (image[285],filter[4],mul_out[715][10]);
mul_8x8bit m2147 (image[286],filter[5],mul_out[715][11]);
mul_8x8bit m2148 (image[312],filter[6],mul_out[716][9]);
mul_8x8bit m2149 (image[313],filter[7],mul_out[716][10]);
mul_8x8bit m2150 (image[314],filter[8],mul_out[716][11]);

adder_8bit ad238 (mul_out[714][9],mul_out[714][10],mul_out[714][11],mul_out[715][9],mul_out[715][10],mul_out[715][11],mul_out[716][9],mul_out[716][10],mul_out[716][11],conv_out[238]);



mul_8x8bit m2151 (image[257],filter[0],mul_out[717][9]);
mul_8x8bit m2152 (image[258],filter[1],mul_out[717][10]);
mul_8x8bit m2153 (image[259],filter[2],mul_out[717][11]);
mul_8x8bit m2154 (image[285],filter[3],mul_out[718][9]);
mul_8x8bit m2155 (image[286],filter[4],mul_out[718][10]);
mul_8x8bit m2156 (image[287],filter[5],mul_out[718][11]);
mul_8x8bit m2157 (image[313],filter[6],mul_out[719][9]);
mul_8x8bit m2158 (image[314],filter[7],mul_out[719][10]);
mul_8x8bit m2159 (image[315],filter[8],mul_out[719][11]);

adder_8bit ad239 (mul_out[717][9],mul_out[717][10],mul_out[717][11],mul_out[718][9],mul_out[718][10],mul_out[718][11],mul_out[719][9],mul_out[719][10],mul_out[719][11],conv_out[239]);



mul_8x8bit m2160 (image[258],filter[0],mul_out[720][9]);
mul_8x8bit m2161 (image[259],filter[1],mul_out[720][10]);
mul_8x8bit m2162 (image[260],filter[2],mul_out[720][11]);
mul_8x8bit m2163 (image[286],filter[3],mul_out[721][9]);
mul_8x8bit m2164 (image[287],filter[4],mul_out[721][10]);
mul_8x8bit m2165 (image[288],filter[5],mul_out[721][11]);
mul_8x8bit m2166 (image[314],filter[6],mul_out[722][9]);
mul_8x8bit m2167 (image[315],filter[7],mul_out[722][10]);
mul_8x8bit m2168 (image[316],filter[8],mul_out[722][11]);

adder_8bit ad240 (mul_out[720][9],mul_out[720][10],mul_out[720][11],mul_out[721][9],mul_out[721][10],mul_out[721][11],mul_out[722][9],mul_out[722][10],mul_out[722][11],conv_out[240]);



mul_8x8bit m2169 (image[259],filter[0],mul_out[723][9]);
mul_8x8bit m2170 (image[260],filter[1],mul_out[723][10]);
mul_8x8bit m2171 (image[261],filter[2],mul_out[723][11]);
mul_8x8bit m2172 (image[287],filter[3],mul_out[724][9]);
mul_8x8bit m2173 (image[288],filter[4],mul_out[724][10]);
mul_8x8bit m2174 (image[289],filter[5],mul_out[724][11]);
mul_8x8bit m2175 (image[315],filter[6],mul_out[725][9]);
mul_8x8bit m2176 (image[316],filter[7],mul_out[725][10]);
mul_8x8bit m2177 (image[317],filter[8],mul_out[725][11]);

adder_8bit ad241 (mul_out[723][9],mul_out[723][10],mul_out[723][11],mul_out[724][9],mul_out[724][10],mul_out[724][11],mul_out[725][9],mul_out[725][10],mul_out[725][11],conv_out[241]);



mul_8x8bit m2178 (image[260],filter[0],mul_out[726][9]);
mul_8x8bit m2179 (image[261],filter[1],mul_out[726][10]);
mul_8x8bit m2180 (image[262],filter[2],mul_out[726][11]);
mul_8x8bit m2181 (image[288],filter[3],mul_out[727][9]);
mul_8x8bit m2182 (image[289],filter[4],mul_out[727][10]);
mul_8x8bit m2183 (image[290],filter[5],mul_out[727][11]);
mul_8x8bit m2184 (image[316],filter[6],mul_out[728][9]);
mul_8x8bit m2185 (image[317],filter[7],mul_out[728][10]);
mul_8x8bit m2186 (image[318],filter[8],mul_out[728][11]);

adder_8bit ad242 (mul_out[726][9],mul_out[726][10],mul_out[726][11],mul_out[727][9],mul_out[727][10],mul_out[727][11],mul_out[728][9],mul_out[728][10],mul_out[728][11],conv_out[242]);



mul_8x8bit m2187 (image[261],filter[0],mul_out[729][9]);
mul_8x8bit m2188 (image[262],filter[1],mul_out[729][10]);
mul_8x8bit m2189 (image[263],filter[2],mul_out[729][11]);
mul_8x8bit m2190 (image[289],filter[3],mul_out[730][9]);
mul_8x8bit m2191 (image[290],filter[4],mul_out[730][10]);
mul_8x8bit m2192 (image[291],filter[5],mul_out[730][11]);
mul_8x8bit m2193 (image[317],filter[6],mul_out[731][9]);
mul_8x8bit m2194 (image[318],filter[7],mul_out[731][10]);
mul_8x8bit m2195 (image[319],filter[8],mul_out[731][11]);

adder_8bit ad243 (mul_out[729][9],mul_out[729][10],mul_out[729][11],mul_out[730][9],mul_out[730][10],mul_out[730][11],mul_out[731][9],mul_out[731][10],mul_out[731][11],conv_out[243]);



mul_8x8bit m2196 (image[262],filter[0],mul_out[732][9]);
mul_8x8bit m2197 (image[263],filter[1],mul_out[732][10]);
mul_8x8bit m2198 (image[264],filter[2],mul_out[732][11]);
mul_8x8bit m2199 (image[290],filter[3],mul_out[733][9]);
mul_8x8bit m2200 (image[291],filter[4],mul_out[733][10]);
mul_8x8bit m2201 (image[292],filter[5],mul_out[733][11]);
mul_8x8bit m2202 (image[318],filter[6],mul_out[734][9]);
mul_8x8bit m2203 (image[319],filter[7],mul_out[734][10]);
mul_8x8bit m2204 (image[320],filter[8],mul_out[734][11]);

adder_8bit ad244 (mul_out[732][9],mul_out[732][10],mul_out[732][11],mul_out[733][9],mul_out[733][10],mul_out[733][11],mul_out[734][9],mul_out[734][10],mul_out[734][11],conv_out[244]);



mul_8x8bit m2205 (image[263],filter[0],mul_out[735][9]);
mul_8x8bit m2206 (image[264],filter[1],mul_out[735][10]);
mul_8x8bit m2207 (image[265],filter[2],mul_out[735][11]);
mul_8x8bit m2208 (image[291],filter[3],mul_out[736][9]);
mul_8x8bit m2209 (image[292],filter[4],mul_out[736][10]);
mul_8x8bit m2210 (image[293],filter[5],mul_out[736][11]);
mul_8x8bit m2211 (image[319],filter[6],mul_out[737][9]);
mul_8x8bit m2212 (image[320],filter[7],mul_out[737][10]);
mul_8x8bit m2213 (image[321],filter[8],mul_out[737][11]);

adder_8bit ad245 (mul_out[735][9],mul_out[735][10],mul_out[735][11],mul_out[736][9],mul_out[736][10],mul_out[736][11],mul_out[737][9],mul_out[737][10],mul_out[737][11],conv_out[245]);



mul_8x8bit m2214 (image[264],filter[0],mul_out[738][9]);
mul_8x8bit m2215 (image[265],filter[1],mul_out[738][10]);
mul_8x8bit m2216 (image[266],filter[2],mul_out[738][11]);
mul_8x8bit m2217 (image[292],filter[3],mul_out[739][9]);
mul_8x8bit m2218 (image[293],filter[4],mul_out[739][10]);
mul_8x8bit m2219 (image[294],filter[5],mul_out[739][11]);
mul_8x8bit m2220 (image[320],filter[6],mul_out[740][9]);
mul_8x8bit m2221 (image[321],filter[7],mul_out[740][10]);
mul_8x8bit m2222 (image[322],filter[8],mul_out[740][11]);

adder_8bit ad246 (mul_out[738][9],mul_out[738][10],mul_out[738][11],mul_out[739][9],mul_out[739][10],mul_out[739][11],mul_out[740][9],mul_out[740][10],mul_out[740][11],conv_out[246]);



mul_8x8bit m2223 (image[265],filter[0],mul_out[741][9]);
mul_8x8bit m2224 (image[266],filter[1],mul_out[741][10]);
mul_8x8bit m2225 (image[267],filter[2],mul_out[741][11]);
mul_8x8bit m2226 (image[293],filter[3],mul_out[742][9]);
mul_8x8bit m2227 (image[294],filter[4],mul_out[742][10]);
mul_8x8bit m2228 (image[295],filter[5],mul_out[742][11]);
mul_8x8bit m2229 (image[321],filter[6],mul_out[743][9]);
mul_8x8bit m2230 (image[322],filter[7],mul_out[743][10]);
mul_8x8bit m2231 (image[323],filter[8],mul_out[743][11]);

adder_8bit ad247 (mul_out[741][9],mul_out[741][10],mul_out[741][11],mul_out[742][9],mul_out[742][10],mul_out[742][11],mul_out[743][9],mul_out[743][10],mul_out[743][11],conv_out[247]);



mul_8x8bit m2232 (image[266],filter[0],mul_out[744][9]);
mul_8x8bit m2233 (image[267],filter[1],mul_out[744][10]);
mul_8x8bit m2234 (image[268],filter[2],mul_out[744][11]);
mul_8x8bit m2235 (image[294],filter[3],mul_out[745][9]);
mul_8x8bit m2236 (image[295],filter[4],mul_out[745][10]);
mul_8x8bit m2237 (image[296],filter[5],mul_out[745][11]);
mul_8x8bit m2238 (image[322],filter[6],mul_out[746][9]);
mul_8x8bit m2239 (image[323],filter[7],mul_out[746][10]);
mul_8x8bit m2240 (image[324],filter[8],mul_out[746][11]);

adder_8bit ad248 (mul_out[744][9],mul_out[744][10],mul_out[744][11],mul_out[745][9],mul_out[745][10],mul_out[745][11],mul_out[746][9],mul_out[746][10],mul_out[746][11],conv_out[248]);



mul_8x8bit m2241 (image[267],filter[0],mul_out[747][9]);
mul_8x8bit m2242 (image[268],filter[1],mul_out[747][10]);
mul_8x8bit m2243 (image[269],filter[2],mul_out[747][11]);
mul_8x8bit m2244 (image[295],filter[3],mul_out[748][9]);
mul_8x8bit m2245 (image[296],filter[4],mul_out[748][10]);
mul_8x8bit m2246 (image[297],filter[5],mul_out[748][11]);
mul_8x8bit m2247 (image[323],filter[6],mul_out[749][9]);
mul_8x8bit m2248 (image[324],filter[7],mul_out[749][10]);
mul_8x8bit m2249 (image[325],filter[8],mul_out[749][11]);

adder_8bit ad249 (mul_out[747][9],mul_out[747][10],mul_out[747][11],mul_out[748][9],mul_out[748][10],mul_out[748][11],mul_out[749][9],mul_out[749][10],mul_out[749][11],conv_out[249]);



mul_8x8bit m2250 (image[268],filter[0],mul_out[750][9]);
mul_8x8bit m2251 (image[269],filter[1],mul_out[750][10]);
mul_8x8bit m2252 (image[270],filter[2],mul_out[750][11]);
mul_8x8bit m2253 (image[296],filter[3],mul_out[751][9]);
mul_8x8bit m2254 (image[297],filter[4],mul_out[751][10]);
mul_8x8bit m2255 (image[298],filter[5],mul_out[751][11]);
mul_8x8bit m2256 (image[324],filter[6],mul_out[752][9]);
mul_8x8bit m2257 (image[325],filter[7],mul_out[752][10]);
mul_8x8bit m2258 (image[326],filter[8],mul_out[752][11]);

adder_8bit ad250 (mul_out[750][9],mul_out[750][10],mul_out[750][11],mul_out[751][9],mul_out[751][10],mul_out[751][11],mul_out[752][9],mul_out[752][10],mul_out[752][11],conv_out[250]);



mul_8x8bit m2259 (image[269],filter[0],mul_out[753][9]);
mul_8x8bit m2260 (image[270],filter[1],mul_out[753][10]);
mul_8x8bit m2261 (image[271],filter[2],mul_out[753][11]);
mul_8x8bit m2262 (image[297],filter[3],mul_out[754][9]);
mul_8x8bit m2263 (image[298],filter[4],mul_out[754][10]);
mul_8x8bit m2264 (image[299],filter[5],mul_out[754][11]);
mul_8x8bit m2265 (image[325],filter[6],mul_out[755][9]);
mul_8x8bit m2266 (image[326],filter[7],mul_out[755][10]);
mul_8x8bit m2267 (image[327],filter[8],mul_out[755][11]);

adder_8bit ad251 (mul_out[753][9],mul_out[753][10],mul_out[753][11],mul_out[754][9],mul_out[754][10],mul_out[754][11],mul_out[755][9],mul_out[755][10],mul_out[755][11],conv_out[251]);



mul_8x8bit m2268 (image[270],filter[0],mul_out[756][9]);
mul_8x8bit m2269 (image[271],filter[1],mul_out[756][10]);
mul_8x8bit m2270 (image[272],filter[2],mul_out[756][11]);
mul_8x8bit m2271 (image[298],filter[3],mul_out[757][9]);
mul_8x8bit m2272 (image[299],filter[4],mul_out[757][10]);
mul_8x8bit m2273 (image[300],filter[5],mul_out[757][11]);
mul_8x8bit m2274 (image[326],filter[6],mul_out[758][9]);
mul_8x8bit m2275 (image[327],filter[7],mul_out[758][10]);
mul_8x8bit m2276 (image[328],filter[8],mul_out[758][11]);

adder_8bit ad252 (mul_out[756][9],mul_out[756][10],mul_out[756][11],mul_out[757][9],mul_out[757][10],mul_out[757][11],mul_out[758][9],mul_out[758][10],mul_out[758][11],conv_out[252]);



mul_8x8bit m2277 (image[271],filter[0],mul_out[759][9]);
mul_8x8bit m2278 (image[272],filter[1],mul_out[759][10]);
mul_8x8bit m2279 (image[273],filter[2],mul_out[759][11]);
mul_8x8bit m2280 (image[299],filter[3],mul_out[760][9]);
mul_8x8bit m2281 (image[300],filter[4],mul_out[760][10]);
mul_8x8bit m2282 (image[301],filter[5],mul_out[760][11]);
mul_8x8bit m2283 (image[327],filter[6],mul_out[761][9]);
mul_8x8bit m2284 (image[328],filter[7],mul_out[761][10]);
mul_8x8bit m2285 (image[329],filter[8],mul_out[761][11]);

adder_8bit ad253 (mul_out[759][9],mul_out[759][10],mul_out[759][11],mul_out[760][9],mul_out[760][10],mul_out[760][11],mul_out[761][9],mul_out[761][10],mul_out[761][11],conv_out[253]);



mul_8x8bit m2286 (image[272],filter[0],mul_out[762][9]);
mul_8x8bit m2287 (image[273],filter[1],mul_out[762][10]);
mul_8x8bit m2288 (image[274],filter[2],mul_out[762][11]);
mul_8x8bit m2289 (image[300],filter[3],mul_out[763][9]);
mul_8x8bit m2290 (image[301],filter[4],mul_out[763][10]);
mul_8x8bit m2291 (image[302],filter[5],mul_out[763][11]);
mul_8x8bit m2292 (image[328],filter[6],mul_out[764][9]);
mul_8x8bit m2293 (image[329],filter[7],mul_out[764][10]);
mul_8x8bit m2294 (image[330],filter[8],mul_out[764][11]);

adder_8bit ad254 (mul_out[762][9],mul_out[762][10],mul_out[762][11],mul_out[763][9],mul_out[763][10],mul_out[763][11],mul_out[764][9],mul_out[764][10],mul_out[764][11],conv_out[254]);



mul_8x8bit m2295 (image[273],filter[0],mul_out[765][9]);
mul_8x8bit m2296 (image[274],filter[1],mul_out[765][10]);
mul_8x8bit m2297 (image[275],filter[2],mul_out[765][11]);
mul_8x8bit m2298 (image[301],filter[3],mul_out[766][9]);
mul_8x8bit m2299 (image[302],filter[4],mul_out[766][10]);
mul_8x8bit m2300 (image[303],filter[5],mul_out[766][11]);
mul_8x8bit m2301 (image[329],filter[6],mul_out[767][9]);
mul_8x8bit m2302 (image[330],filter[7],mul_out[767][10]);
mul_8x8bit m2303 (image[331],filter[8],mul_out[767][11]);

adder_8bit ad255 (mul_out[765][9],mul_out[765][10],mul_out[765][11],mul_out[766][9],mul_out[766][10],mul_out[766][11],mul_out[767][9],mul_out[767][10],mul_out[767][11],conv_out[255]);



mul_8x8bit m2304 (image[274],filter[0],mul_out[768][9]);
mul_8x8bit m2305 (image[275],filter[1],mul_out[768][10]);
mul_8x8bit m2306 (image[276],filter[2],mul_out[768][11]);
mul_8x8bit m2307 (image[302],filter[3],mul_out[769][9]);
mul_8x8bit m2308 (image[303],filter[4],mul_out[769][10]);
mul_8x8bit m2309 (image[304],filter[5],mul_out[769][11]);
mul_8x8bit m2310 (image[330],filter[6],mul_out[770][9]);
mul_8x8bit m2311 (image[331],filter[7],mul_out[770][10]);
mul_8x8bit m2312 (image[332],filter[8],mul_out[770][11]);

adder_8bit ad256 (mul_out[768][9],mul_out[768][10],mul_out[768][11],mul_out[769][9],mul_out[769][10],mul_out[769][11],mul_out[770][9],mul_out[770][10],mul_out[770][11],conv_out[256]);



mul_8x8bit m2313 (image[275],filter[0],mul_out[771][9]);
mul_8x8bit m2314 (image[276],filter[1],mul_out[771][10]);
mul_8x8bit m2315 (image[277],filter[2],mul_out[771][11]);
mul_8x8bit m2316 (image[303],filter[3],mul_out[772][9]);
mul_8x8bit m2317 (image[304],filter[4],mul_out[772][10]);
mul_8x8bit m2318 (image[305],filter[5],mul_out[772][11]);
mul_8x8bit m2319 (image[331],filter[6],mul_out[773][9]);
mul_8x8bit m2320 (image[332],filter[7],mul_out[773][10]);
mul_8x8bit m2321 (image[333],filter[8],mul_out[773][11]);

adder_8bit ad257 (mul_out[771][9],mul_out[771][10],mul_out[771][11],mul_out[772][9],mul_out[772][10],mul_out[772][11],mul_out[773][9],mul_out[773][10],mul_out[773][11],conv_out[257]);



mul_8x8bit m2322 (image[276],filter[0],mul_out[774][9]);
mul_8x8bit m2323 (image[277],filter[1],mul_out[774][10]);
mul_8x8bit m2324 (image[278],filter[2],mul_out[774][11]);
mul_8x8bit m2325 (image[304],filter[3],mul_out[775][9]);
mul_8x8bit m2326 (image[305],filter[4],mul_out[775][10]);
mul_8x8bit m2327 (image[306],filter[5],mul_out[775][11]);
mul_8x8bit m2328 (image[332],filter[6],mul_out[776][9]);
mul_8x8bit m2329 (image[333],filter[7],mul_out[776][10]);
mul_8x8bit m2330 (image[334],filter[8],mul_out[776][11]);

adder_8bit ad258 (mul_out[774][9],mul_out[774][10],mul_out[774][11],mul_out[775][9],mul_out[775][10],mul_out[775][11],mul_out[776][9],mul_out[776][10],mul_out[776][11],conv_out[258]);



mul_8x8bit m2331 (image[277],filter[0],mul_out[777][9]);
mul_8x8bit m2332 (image[278],filter[1],mul_out[777][10]);
mul_8x8bit m2333 (image[279],filter[2],mul_out[777][11]);
mul_8x8bit m2334 (image[305],filter[3],mul_out[778][9]);
mul_8x8bit m2335 (image[306],filter[4],mul_out[778][10]);
mul_8x8bit m2336 (image[307],filter[5],mul_out[778][11]);
mul_8x8bit m2337 (image[333],filter[6],mul_out[779][9]);
mul_8x8bit m2338 (image[334],filter[7],mul_out[779][10]);
mul_8x8bit m2339 (image[335],filter[8],mul_out[779][11]);

adder_8bit ad259 (mul_out[777][9],mul_out[777][10],mul_out[777][11],mul_out[778][9],mul_out[778][10],mul_out[778][11],mul_out[779][9],mul_out[779][10],mul_out[779][11],conv_out[259]);



mul_8x8bit m2340 (image[280],filter[0],mul_out[780][10]);
mul_8x8bit m2341 (image[281],filter[1],mul_out[780][11]);
mul_8x8bit m2342 (image[282],filter[2],mul_out[780][12]);
mul_8x8bit m2343 (image[308],filter[3],mul_out[781][10]);
mul_8x8bit m2344 (image[309],filter[4],mul_out[781][11]);
mul_8x8bit m2345 (image[310],filter[5],mul_out[781][12]);
mul_8x8bit m2346 (image[336],filter[6],mul_out[782][10]);
mul_8x8bit m2347 (image[337],filter[7],mul_out[782][11]);
mul_8x8bit m2348 (image[338],filter[8],mul_out[782][12]);

adder_8bit ad260 (mul_out[780][10],mul_out[780][11],mul_out[780][12],mul_out[781][10],mul_out[781][11],mul_out[781][12],mul_out[782][10],mul_out[782][11],mul_out[782][12],conv_out[260]);



mul_8x8bit m2349 (image[281],filter[0],mul_out[783][10]);
mul_8x8bit m2350 (image[282],filter[1],mul_out[783][11]);
mul_8x8bit m2351 (image[283],filter[2],mul_out[783][12]);
mul_8x8bit m2352 (image[309],filter[3],mul_out[784][10]);
mul_8x8bit m2353 (image[310],filter[4],mul_out[784][11]);
mul_8x8bit m2354 (image[311],filter[5],mul_out[784][12]);
mul_8x8bit m2355 (image[337],filter[6],mul_out[785][10]);
mul_8x8bit m2356 (image[338],filter[7],mul_out[785][11]);
mul_8x8bit m2357 (image[339],filter[8],mul_out[785][12]);

adder_8bit ad261 (mul_out[783][10],mul_out[783][11],mul_out[783][12],mul_out[784][10],mul_out[784][11],mul_out[784][12],mul_out[785][10],mul_out[785][11],mul_out[785][12],conv_out[261]);



mul_8x8bit m2358 (image[282],filter[0],mul_out[786][10]);
mul_8x8bit m2359 (image[283],filter[1],mul_out[786][11]);
mul_8x8bit m2360 (image[284],filter[2],mul_out[786][12]);
mul_8x8bit m2361 (image[310],filter[3],mul_out[787][10]);
mul_8x8bit m2362 (image[311],filter[4],mul_out[787][11]);
mul_8x8bit m2363 (image[312],filter[5],mul_out[787][12]);
mul_8x8bit m2364 (image[338],filter[6],mul_out[788][10]);
mul_8x8bit m2365 (image[339],filter[7],mul_out[788][11]);
mul_8x8bit m2366 (image[340],filter[8],mul_out[788][12]);

adder_8bit ad262 (mul_out[786][10],mul_out[786][11],mul_out[786][12],mul_out[787][10],mul_out[787][11],mul_out[787][12],mul_out[788][10],mul_out[788][11],mul_out[788][12],conv_out[262]);



mul_8x8bit m2367 (image[283],filter[0],mul_out[789][10]);
mul_8x8bit m2368 (image[284],filter[1],mul_out[789][11]);
mul_8x8bit m2369 (image[285],filter[2],mul_out[789][12]);
mul_8x8bit m2370 (image[311],filter[3],mul_out[790][10]);
mul_8x8bit m2371 (image[312],filter[4],mul_out[790][11]);
mul_8x8bit m2372 (image[313],filter[5],mul_out[790][12]);
mul_8x8bit m2373 (image[339],filter[6],mul_out[791][10]);
mul_8x8bit m2374 (image[340],filter[7],mul_out[791][11]);
mul_8x8bit m2375 (image[341],filter[8],mul_out[791][12]);

adder_8bit ad263 (mul_out[789][10],mul_out[789][11],mul_out[789][12],mul_out[790][10],mul_out[790][11],mul_out[790][12],mul_out[791][10],mul_out[791][11],mul_out[791][12],conv_out[263]);



mul_8x8bit m2376 (image[284],filter[0],mul_out[792][10]);
mul_8x8bit m2377 (image[285],filter[1],mul_out[792][11]);
mul_8x8bit m2378 (image[286],filter[2],mul_out[792][12]);
mul_8x8bit m2379 (image[312],filter[3],mul_out[793][10]);
mul_8x8bit m2380 (image[313],filter[4],mul_out[793][11]);
mul_8x8bit m2381 (image[314],filter[5],mul_out[793][12]);
mul_8x8bit m2382 (image[340],filter[6],mul_out[794][10]);
mul_8x8bit m2383 (image[341],filter[7],mul_out[794][11]);
mul_8x8bit m2384 (image[342],filter[8],mul_out[794][12]);

adder_8bit ad264 (mul_out[792][10],mul_out[792][11],mul_out[792][12],mul_out[793][10],mul_out[793][11],mul_out[793][12],mul_out[794][10],mul_out[794][11],mul_out[794][12],conv_out[264]);



mul_8x8bit m2385 (image[285],filter[0],mul_out[795][10]);
mul_8x8bit m2386 (image[286],filter[1],mul_out[795][11]);
mul_8x8bit m2387 (image[287],filter[2],mul_out[795][12]);
mul_8x8bit m2388 (image[313],filter[3],mul_out[796][10]);
mul_8x8bit m2389 (image[314],filter[4],mul_out[796][11]);
mul_8x8bit m2390 (image[315],filter[5],mul_out[796][12]);
mul_8x8bit m2391 (image[341],filter[6],mul_out[797][10]);
mul_8x8bit m2392 (image[342],filter[7],mul_out[797][11]);
mul_8x8bit m2393 (image[343],filter[8],mul_out[797][12]);

adder_8bit ad265 (mul_out[795][10],mul_out[795][11],mul_out[795][12],mul_out[796][10],mul_out[796][11],mul_out[796][12],mul_out[797][10],mul_out[797][11],mul_out[797][12],conv_out[265]);



mul_8x8bit m2394 (image[286],filter[0],mul_out[798][10]);
mul_8x8bit m2395 (image[287],filter[1],mul_out[798][11]);
mul_8x8bit m2396 (image[288],filter[2],mul_out[798][12]);
mul_8x8bit m2397 (image[314],filter[3],mul_out[799][10]);
mul_8x8bit m2398 (image[315],filter[4],mul_out[799][11]);
mul_8x8bit m2399 (image[316],filter[5],mul_out[799][12]);
mul_8x8bit m2400 (image[342],filter[6],mul_out[800][10]);
mul_8x8bit m2401 (image[343],filter[7],mul_out[800][11]);
mul_8x8bit m2402 (image[344],filter[8],mul_out[800][12]);

adder_8bit ad266 (mul_out[798][10],mul_out[798][11],mul_out[798][12],mul_out[799][10],mul_out[799][11],mul_out[799][12],mul_out[800][10],mul_out[800][11],mul_out[800][12],conv_out[266]);



mul_8x8bit m2403 (image[287],filter[0],mul_out[801][10]);
mul_8x8bit m2404 (image[288],filter[1],mul_out[801][11]);
mul_8x8bit m2405 (image[289],filter[2],mul_out[801][12]);
mul_8x8bit m2406 (image[315],filter[3],mul_out[802][10]);
mul_8x8bit m2407 (image[316],filter[4],mul_out[802][11]);
mul_8x8bit m2408 (image[317],filter[5],mul_out[802][12]);
mul_8x8bit m2409 (image[343],filter[6],mul_out[803][10]);
mul_8x8bit m2410 (image[344],filter[7],mul_out[803][11]);
mul_8x8bit m2411 (image[345],filter[8],mul_out[803][12]);

adder_8bit ad267 (mul_out[801][10],mul_out[801][11],mul_out[801][12],mul_out[802][10],mul_out[802][11],mul_out[802][12],mul_out[803][10],mul_out[803][11],mul_out[803][12],conv_out[267]);



mul_8x8bit m2412 (image[288],filter[0],mul_out[804][10]);
mul_8x8bit m2413 (image[289],filter[1],mul_out[804][11]);
mul_8x8bit m2414 (image[290],filter[2],mul_out[804][12]);
mul_8x8bit m2415 (image[316],filter[3],mul_out[805][10]);
mul_8x8bit m2416 (image[317],filter[4],mul_out[805][11]);
mul_8x8bit m2417 (image[318],filter[5],mul_out[805][12]);
mul_8x8bit m2418 (image[344],filter[6],mul_out[806][10]);
mul_8x8bit m2419 (image[345],filter[7],mul_out[806][11]);
mul_8x8bit m2420 (image[346],filter[8],mul_out[806][12]);

adder_8bit ad268 (mul_out[804][10],mul_out[804][11],mul_out[804][12],mul_out[805][10],mul_out[805][11],mul_out[805][12],mul_out[806][10],mul_out[806][11],mul_out[806][12],conv_out[268]);



mul_8x8bit m2421 (image[289],filter[0],mul_out[807][10]);
mul_8x8bit m2422 (image[290],filter[1],mul_out[807][11]);
mul_8x8bit m2423 (image[291],filter[2],mul_out[807][12]);
mul_8x8bit m2424 (image[317],filter[3],mul_out[808][10]);
mul_8x8bit m2425 (image[318],filter[4],mul_out[808][11]);
mul_8x8bit m2426 (image[319],filter[5],mul_out[808][12]);
mul_8x8bit m2427 (image[345],filter[6],mul_out[809][10]);
mul_8x8bit m2428 (image[346],filter[7],mul_out[809][11]);
mul_8x8bit m2429 (image[347],filter[8],mul_out[809][12]);

adder_8bit ad269 (mul_out[807][10],mul_out[807][11],mul_out[807][12],mul_out[808][10],mul_out[808][11],mul_out[808][12],mul_out[809][10],mul_out[809][11],mul_out[809][12],conv_out[269]);



mul_8x8bit m2430 (image[290],filter[0],mul_out[810][10]);
mul_8x8bit m2431 (image[291],filter[1],mul_out[810][11]);
mul_8x8bit m2432 (image[292],filter[2],mul_out[810][12]);
mul_8x8bit m2433 (image[318],filter[3],mul_out[811][10]);
mul_8x8bit m2434 (image[319],filter[4],mul_out[811][11]);
mul_8x8bit m2435 (image[320],filter[5],mul_out[811][12]);
mul_8x8bit m2436 (image[346],filter[6],mul_out[812][10]);
mul_8x8bit m2437 (image[347],filter[7],mul_out[812][11]);
mul_8x8bit m2438 (image[348],filter[8],mul_out[812][12]);

adder_8bit ad270 (mul_out[810][10],mul_out[810][11],mul_out[810][12],mul_out[811][10],mul_out[811][11],mul_out[811][12],mul_out[812][10],mul_out[812][11],mul_out[812][12],conv_out[270]);



mul_8x8bit m2439 (image[291],filter[0],mul_out[813][10]);
mul_8x8bit m2440 (image[292],filter[1],mul_out[813][11]);
mul_8x8bit m2441 (image[293],filter[2],mul_out[813][12]);
mul_8x8bit m2442 (image[319],filter[3],mul_out[814][10]);
mul_8x8bit m2443 (image[320],filter[4],mul_out[814][11]);
mul_8x8bit m2444 (image[321],filter[5],mul_out[814][12]);
mul_8x8bit m2445 (image[347],filter[6],mul_out[815][10]);
mul_8x8bit m2446 (image[348],filter[7],mul_out[815][11]);
mul_8x8bit m2447 (image[349],filter[8],mul_out[815][12]);

adder_8bit ad271 (mul_out[813][10],mul_out[813][11],mul_out[813][12],mul_out[814][10],mul_out[814][11],mul_out[814][12],mul_out[815][10],mul_out[815][11],mul_out[815][12],conv_out[271]);



mul_8x8bit m2448 (image[292],filter[0],mul_out[816][10]);
mul_8x8bit m2449 (image[293],filter[1],mul_out[816][11]);
mul_8x8bit m2450 (image[294],filter[2],mul_out[816][12]);
mul_8x8bit m2451 (image[320],filter[3],mul_out[817][10]);
mul_8x8bit m2452 (image[321],filter[4],mul_out[817][11]);
mul_8x8bit m2453 (image[322],filter[5],mul_out[817][12]);
mul_8x8bit m2454 (image[348],filter[6],mul_out[818][10]);
mul_8x8bit m2455 (image[349],filter[7],mul_out[818][11]);
mul_8x8bit m2456 (image[350],filter[8],mul_out[818][12]);

adder_8bit ad272 (mul_out[816][10],mul_out[816][11],mul_out[816][12],mul_out[817][10],mul_out[817][11],mul_out[817][12],mul_out[818][10],mul_out[818][11],mul_out[818][12],conv_out[272]);



mul_8x8bit m2457 (image[293],filter[0],mul_out[819][10]);
mul_8x8bit m2458 (image[294],filter[1],mul_out[819][11]);
mul_8x8bit m2459 (image[295],filter[2],mul_out[819][12]);
mul_8x8bit m2460 (image[321],filter[3],mul_out[820][10]);
mul_8x8bit m2461 (image[322],filter[4],mul_out[820][11]);
mul_8x8bit m2462 (image[323],filter[5],mul_out[820][12]);
mul_8x8bit m2463 (image[349],filter[6],mul_out[821][10]);
mul_8x8bit m2464 (image[350],filter[7],mul_out[821][11]);
mul_8x8bit m2465 (image[351],filter[8],mul_out[821][12]);

adder_8bit ad273 (mul_out[819][10],mul_out[819][11],mul_out[819][12],mul_out[820][10],mul_out[820][11],mul_out[820][12],mul_out[821][10],mul_out[821][11],mul_out[821][12],conv_out[273]);



mul_8x8bit m2466 (image[294],filter[0],mul_out[822][10]);
mul_8x8bit m2467 (image[295],filter[1],mul_out[822][11]);
mul_8x8bit m2468 (image[296],filter[2],mul_out[822][12]);
mul_8x8bit m2469 (image[322],filter[3],mul_out[823][10]);
mul_8x8bit m2470 (image[323],filter[4],mul_out[823][11]);
mul_8x8bit m2471 (image[324],filter[5],mul_out[823][12]);
mul_8x8bit m2472 (image[350],filter[6],mul_out[824][10]);
mul_8x8bit m2473 (image[351],filter[7],mul_out[824][11]);
mul_8x8bit m2474 (image[352],filter[8],mul_out[824][12]);

adder_8bit ad274 (mul_out[822][10],mul_out[822][11],mul_out[822][12],mul_out[823][10],mul_out[823][11],mul_out[823][12],mul_out[824][10],mul_out[824][11],mul_out[824][12],conv_out[274]);



mul_8x8bit m2475 (image[295],filter[0],mul_out[825][10]);
mul_8x8bit m2476 (image[296],filter[1],mul_out[825][11]);
mul_8x8bit m2477 (image[297],filter[2],mul_out[825][12]);
mul_8x8bit m2478 (image[323],filter[3],mul_out[826][10]);
mul_8x8bit m2479 (image[324],filter[4],mul_out[826][11]);
mul_8x8bit m2480 (image[325],filter[5],mul_out[826][12]);
mul_8x8bit m2481 (image[351],filter[6],mul_out[827][10]);
mul_8x8bit m2482 (image[352],filter[7],mul_out[827][11]);
mul_8x8bit m2483 (image[353],filter[8],mul_out[827][12]);

adder_8bit ad275 (mul_out[825][10],mul_out[825][11],mul_out[825][12],mul_out[826][10],mul_out[826][11],mul_out[826][12],mul_out[827][10],mul_out[827][11],mul_out[827][12],conv_out[275]);



mul_8x8bit m2484 (image[296],filter[0],mul_out[828][10]);
mul_8x8bit m2485 (image[297],filter[1],mul_out[828][11]);
mul_8x8bit m2486 (image[298],filter[2],mul_out[828][12]);
mul_8x8bit m2487 (image[324],filter[3],mul_out[829][10]);
mul_8x8bit m2488 (image[325],filter[4],mul_out[829][11]);
mul_8x8bit m2489 (image[326],filter[5],mul_out[829][12]);
mul_8x8bit m2490 (image[352],filter[6],mul_out[830][10]);
mul_8x8bit m2491 (image[353],filter[7],mul_out[830][11]);
mul_8x8bit m2492 (image[354],filter[8],mul_out[830][12]);

adder_8bit ad276 (mul_out[828][10],mul_out[828][11],mul_out[828][12],mul_out[829][10],mul_out[829][11],mul_out[829][12],mul_out[830][10],mul_out[830][11],mul_out[830][12],conv_out[276]);



mul_8x8bit m2493 (image[297],filter[0],mul_out[831][10]);
mul_8x8bit m2494 (image[298],filter[1],mul_out[831][11]);
mul_8x8bit m2495 (image[299],filter[2],mul_out[831][12]);
mul_8x8bit m2496 (image[325],filter[3],mul_out[832][10]);
mul_8x8bit m2497 (image[326],filter[4],mul_out[832][11]);
mul_8x8bit m2498 (image[327],filter[5],mul_out[832][12]);
mul_8x8bit m2499 (image[353],filter[6],mul_out[833][10]);
mul_8x8bit m2500 (image[354],filter[7],mul_out[833][11]);
mul_8x8bit m2501 (image[355],filter[8],mul_out[833][12]);

adder_8bit ad277 (mul_out[831][10],mul_out[831][11],mul_out[831][12],mul_out[832][10],mul_out[832][11],mul_out[832][12],mul_out[833][10],mul_out[833][11],mul_out[833][12],conv_out[277]);



mul_8x8bit m2502 (image[298],filter[0],mul_out[834][10]);
mul_8x8bit m2503 (image[299],filter[1],mul_out[834][11]);
mul_8x8bit m2504 (image[300],filter[2],mul_out[834][12]);
mul_8x8bit m2505 (image[326],filter[3],mul_out[835][10]);
mul_8x8bit m2506 (image[327],filter[4],mul_out[835][11]);
mul_8x8bit m2507 (image[328],filter[5],mul_out[835][12]);
mul_8x8bit m2508 (image[354],filter[6],mul_out[836][10]);
mul_8x8bit m2509 (image[355],filter[7],mul_out[836][11]);
mul_8x8bit m2510 (image[356],filter[8],mul_out[836][12]);

adder_8bit ad278 (mul_out[834][10],mul_out[834][11],mul_out[834][12],mul_out[835][10],mul_out[835][11],mul_out[835][12],mul_out[836][10],mul_out[836][11],mul_out[836][12],conv_out[278]);



mul_8x8bit m2511 (image[299],filter[0],mul_out[837][10]);
mul_8x8bit m2512 (image[300],filter[1],mul_out[837][11]);
mul_8x8bit m2513 (image[301],filter[2],mul_out[837][12]);
mul_8x8bit m2514 (image[327],filter[3],mul_out[838][10]);
mul_8x8bit m2515 (image[328],filter[4],mul_out[838][11]);
mul_8x8bit m2516 (image[329],filter[5],mul_out[838][12]);
mul_8x8bit m2517 (image[355],filter[6],mul_out[839][10]);
mul_8x8bit m2518 (image[356],filter[7],mul_out[839][11]);
mul_8x8bit m2519 (image[357],filter[8],mul_out[839][12]);

adder_8bit ad279 (mul_out[837][10],mul_out[837][11],mul_out[837][12],mul_out[838][10],mul_out[838][11],mul_out[838][12],mul_out[839][10],mul_out[839][11],mul_out[839][12],conv_out[279]);



mul_8x8bit m2520 (image[300],filter[0],mul_out[840][10]);
mul_8x8bit m2521 (image[301],filter[1],mul_out[840][11]);
mul_8x8bit m2522 (image[302],filter[2],mul_out[840][12]);
mul_8x8bit m2523 (image[328],filter[3],mul_out[841][10]);
mul_8x8bit m2524 (image[329],filter[4],mul_out[841][11]);
mul_8x8bit m2525 (image[330],filter[5],mul_out[841][12]);
mul_8x8bit m2526 (image[356],filter[6],mul_out[842][10]);
mul_8x8bit m2527 (image[357],filter[7],mul_out[842][11]);
mul_8x8bit m2528 (image[358],filter[8],mul_out[842][12]);

adder_8bit ad280 (mul_out[840][10],mul_out[840][11],mul_out[840][12],mul_out[841][10],mul_out[841][11],mul_out[841][12],mul_out[842][10],mul_out[842][11],mul_out[842][12],conv_out[280]);



mul_8x8bit m2529 (image[301],filter[0],mul_out[843][10]);
mul_8x8bit m2530 (image[302],filter[1],mul_out[843][11]);
mul_8x8bit m2531 (image[303],filter[2],mul_out[843][12]);
mul_8x8bit m2532 (image[329],filter[3],mul_out[844][10]);
mul_8x8bit m2533 (image[330],filter[4],mul_out[844][11]);
mul_8x8bit m2534 (image[331],filter[5],mul_out[844][12]);
mul_8x8bit m2535 (image[357],filter[6],mul_out[845][10]);
mul_8x8bit m2536 (image[358],filter[7],mul_out[845][11]);
mul_8x8bit m2537 (image[359],filter[8],mul_out[845][12]);

adder_8bit ad281 (mul_out[843][10],mul_out[843][11],mul_out[843][12],mul_out[844][10],mul_out[844][11],mul_out[844][12],mul_out[845][10],mul_out[845][11],mul_out[845][12],conv_out[281]);



mul_8x8bit m2538 (image[302],filter[0],mul_out[846][10]);
mul_8x8bit m2539 (image[303],filter[1],mul_out[846][11]);
mul_8x8bit m2540 (image[304],filter[2],mul_out[846][12]);
mul_8x8bit m2541 (image[330],filter[3],mul_out[847][10]);
mul_8x8bit m2542 (image[331],filter[4],mul_out[847][11]);
mul_8x8bit m2543 (image[332],filter[5],mul_out[847][12]);
mul_8x8bit m2544 (image[358],filter[6],mul_out[848][10]);
mul_8x8bit m2545 (image[359],filter[7],mul_out[848][11]);
mul_8x8bit m2546 (image[360],filter[8],mul_out[848][12]);

adder_8bit ad282 (mul_out[846][10],mul_out[846][11],mul_out[846][12],mul_out[847][10],mul_out[847][11],mul_out[847][12],mul_out[848][10],mul_out[848][11],mul_out[848][12],conv_out[282]);



mul_8x8bit m2547 (image[303],filter[0],mul_out[849][10]);
mul_8x8bit m2548 (image[304],filter[1],mul_out[849][11]);
mul_8x8bit m2549 (image[305],filter[2],mul_out[849][12]);
mul_8x8bit m2550 (image[331],filter[3],mul_out[850][10]);
mul_8x8bit m2551 (image[332],filter[4],mul_out[850][11]);
mul_8x8bit m2552 (image[333],filter[5],mul_out[850][12]);
mul_8x8bit m2553 (image[359],filter[6],mul_out[851][10]);
mul_8x8bit m2554 (image[360],filter[7],mul_out[851][11]);
mul_8x8bit m2555 (image[361],filter[8],mul_out[851][12]);

adder_8bit ad283 (mul_out[849][10],mul_out[849][11],mul_out[849][12],mul_out[850][10],mul_out[850][11],mul_out[850][12],mul_out[851][10],mul_out[851][11],mul_out[851][12],conv_out[283]);



mul_8x8bit m2556 (image[304],filter[0],mul_out[852][10]);
mul_8x8bit m2557 (image[305],filter[1],mul_out[852][11]);
mul_8x8bit m2558 (image[306],filter[2],mul_out[852][12]);
mul_8x8bit m2559 (image[332],filter[3],mul_out[853][10]);
mul_8x8bit m2560 (image[333],filter[4],mul_out[853][11]);
mul_8x8bit m2561 (image[334],filter[5],mul_out[853][12]);
mul_8x8bit m2562 (image[360],filter[6],mul_out[854][10]);
mul_8x8bit m2563 (image[361],filter[7],mul_out[854][11]);
mul_8x8bit m2564 (image[362],filter[8],mul_out[854][12]);

adder_8bit ad284 (mul_out[852][10],mul_out[852][11],mul_out[852][12],mul_out[853][10],mul_out[853][11],mul_out[853][12],mul_out[854][10],mul_out[854][11],mul_out[854][12],conv_out[284]);



mul_8x8bit m2565 (image[305],filter[0],mul_out[855][10]);
mul_8x8bit m2566 (image[306],filter[1],mul_out[855][11]);
mul_8x8bit m2567 (image[307],filter[2],mul_out[855][12]);
mul_8x8bit m2568 (image[333],filter[3],mul_out[856][10]);
mul_8x8bit m2569 (image[334],filter[4],mul_out[856][11]);
mul_8x8bit m2570 (image[335],filter[5],mul_out[856][12]);
mul_8x8bit m2571 (image[361],filter[6],mul_out[857][10]);
mul_8x8bit m2572 (image[362],filter[7],mul_out[857][11]);
mul_8x8bit m2573 (image[363],filter[8],mul_out[857][12]);

adder_8bit ad285 (mul_out[855][10],mul_out[855][11],mul_out[855][12],mul_out[856][10],mul_out[856][11],mul_out[856][12],mul_out[857][10],mul_out[857][11],mul_out[857][12],conv_out[285]);



mul_8x8bit m2574 (image[308],filter[0],mul_out[858][11]);
mul_8x8bit m2575 (image[309],filter[1],mul_out[858][12]);
mul_8x8bit m2576 (image[310],filter[2],mul_out[858][13]);
mul_8x8bit m2577 (image[336],filter[3],mul_out[859][11]);
mul_8x8bit m2578 (image[337],filter[4],mul_out[859][12]);
mul_8x8bit m2579 (image[338],filter[5],mul_out[859][13]);
mul_8x8bit m2580 (image[364],filter[6],mul_out[860][11]);
mul_8x8bit m2581 (image[365],filter[7],mul_out[860][12]);
mul_8x8bit m2582 (image[366],filter[8],mul_out[860][13]);

adder_8bit ad286 (mul_out[858][11],mul_out[858][12],mul_out[858][13],mul_out[859][11],mul_out[859][12],mul_out[859][13],mul_out[860][11],mul_out[860][12],mul_out[860][13],conv_out[286]);



mul_8x8bit m2583 (image[309],filter[0],mul_out[861][11]);
mul_8x8bit m2584 (image[310],filter[1],mul_out[861][12]);
mul_8x8bit m2585 (image[311],filter[2],mul_out[861][13]);
mul_8x8bit m2586 (image[337],filter[3],mul_out[862][11]);
mul_8x8bit m2587 (image[338],filter[4],mul_out[862][12]);
mul_8x8bit m2588 (image[339],filter[5],mul_out[862][13]);
mul_8x8bit m2589 (image[365],filter[6],mul_out[863][11]);
mul_8x8bit m2590 (image[366],filter[7],mul_out[863][12]);
mul_8x8bit m2591 (image[367],filter[8],mul_out[863][13]);

adder_8bit ad287 (mul_out[861][11],mul_out[861][12],mul_out[861][13],mul_out[862][11],mul_out[862][12],mul_out[862][13],mul_out[863][11],mul_out[863][12],mul_out[863][13],conv_out[287]);



mul_8x8bit m2592 (image[310],filter[0],mul_out[864][11]);
mul_8x8bit m2593 (image[311],filter[1],mul_out[864][12]);
mul_8x8bit m2594 (image[312],filter[2],mul_out[864][13]);
mul_8x8bit m2595 (image[338],filter[3],mul_out[865][11]);
mul_8x8bit m2596 (image[339],filter[4],mul_out[865][12]);
mul_8x8bit m2597 (image[340],filter[5],mul_out[865][13]);
mul_8x8bit m2598 (image[366],filter[6],mul_out[866][11]);
mul_8x8bit m2599 (image[367],filter[7],mul_out[866][12]);
mul_8x8bit m2600 (image[368],filter[8],mul_out[866][13]);

adder_8bit ad288 (mul_out[864][11],mul_out[864][12],mul_out[864][13],mul_out[865][11],mul_out[865][12],mul_out[865][13],mul_out[866][11],mul_out[866][12],mul_out[866][13],conv_out[288]);



mul_8x8bit m2601 (image[311],filter[0],mul_out[867][11]);
mul_8x8bit m2602 (image[312],filter[1],mul_out[867][12]);
mul_8x8bit m2603 (image[313],filter[2],mul_out[867][13]);
mul_8x8bit m2604 (image[339],filter[3],mul_out[868][11]);
mul_8x8bit m2605 (image[340],filter[4],mul_out[868][12]);
mul_8x8bit m2606 (image[341],filter[5],mul_out[868][13]);
mul_8x8bit m2607 (image[367],filter[6],mul_out[869][11]);
mul_8x8bit m2608 (image[368],filter[7],mul_out[869][12]);
mul_8x8bit m2609 (image[369],filter[8],mul_out[869][13]);

adder_8bit ad289 (mul_out[867][11],mul_out[867][12],mul_out[867][13],mul_out[868][11],mul_out[868][12],mul_out[868][13],mul_out[869][11],mul_out[869][12],mul_out[869][13],conv_out[289]);



mul_8x8bit m2610 (image[312],filter[0],mul_out[870][11]);
mul_8x8bit m2611 (image[313],filter[1],mul_out[870][12]);
mul_8x8bit m2612 (image[314],filter[2],mul_out[870][13]);
mul_8x8bit m2613 (image[340],filter[3],mul_out[871][11]);
mul_8x8bit m2614 (image[341],filter[4],mul_out[871][12]);
mul_8x8bit m2615 (image[342],filter[5],mul_out[871][13]);
mul_8x8bit m2616 (image[368],filter[6],mul_out[872][11]);
mul_8x8bit m2617 (image[369],filter[7],mul_out[872][12]);
mul_8x8bit m2618 (image[370],filter[8],mul_out[872][13]);

adder_8bit ad290 (mul_out[870][11],mul_out[870][12],mul_out[870][13],mul_out[871][11],mul_out[871][12],mul_out[871][13],mul_out[872][11],mul_out[872][12],mul_out[872][13],conv_out[290]);



mul_8x8bit m2619 (image[313],filter[0],mul_out[873][11]);
mul_8x8bit m2620 (image[314],filter[1],mul_out[873][12]);
mul_8x8bit m2621 (image[315],filter[2],mul_out[873][13]);
mul_8x8bit m2622 (image[341],filter[3],mul_out[874][11]);
mul_8x8bit m2623 (image[342],filter[4],mul_out[874][12]);
mul_8x8bit m2624 (image[343],filter[5],mul_out[874][13]);
mul_8x8bit m2625 (image[369],filter[6],mul_out[875][11]);
mul_8x8bit m2626 (image[370],filter[7],mul_out[875][12]);
mul_8x8bit m2627 (image[371],filter[8],mul_out[875][13]);

adder_8bit ad291 (mul_out[873][11],mul_out[873][12],mul_out[873][13],mul_out[874][11],mul_out[874][12],mul_out[874][13],mul_out[875][11],mul_out[875][12],mul_out[875][13],conv_out[291]);



mul_8x8bit m2628 (image[314],filter[0],mul_out[876][11]);
mul_8x8bit m2629 (image[315],filter[1],mul_out[876][12]);
mul_8x8bit m2630 (image[316],filter[2],mul_out[876][13]);
mul_8x8bit m2631 (image[342],filter[3],mul_out[877][11]);
mul_8x8bit m2632 (image[343],filter[4],mul_out[877][12]);
mul_8x8bit m2633 (image[344],filter[5],mul_out[877][13]);
mul_8x8bit m2634 (image[370],filter[6],mul_out[878][11]);
mul_8x8bit m2635 (image[371],filter[7],mul_out[878][12]);
mul_8x8bit m2636 (image[372],filter[8],mul_out[878][13]);

adder_8bit ad292 (mul_out[876][11],mul_out[876][12],mul_out[876][13],mul_out[877][11],mul_out[877][12],mul_out[877][13],mul_out[878][11],mul_out[878][12],mul_out[878][13],conv_out[292]);



mul_8x8bit m2637 (image[315],filter[0],mul_out[879][11]);
mul_8x8bit m2638 (image[316],filter[1],mul_out[879][12]);
mul_8x8bit m2639 (image[317],filter[2],mul_out[879][13]);
mul_8x8bit m2640 (image[343],filter[3],mul_out[880][11]);
mul_8x8bit m2641 (image[344],filter[4],mul_out[880][12]);
mul_8x8bit m2642 (image[345],filter[5],mul_out[880][13]);
mul_8x8bit m2643 (image[371],filter[6],mul_out[881][11]);
mul_8x8bit m2644 (image[372],filter[7],mul_out[881][12]);
mul_8x8bit m2645 (image[373],filter[8],mul_out[881][13]);

adder_8bit ad293 (mul_out[879][11],mul_out[879][12],mul_out[879][13],mul_out[880][11],mul_out[880][12],mul_out[880][13],mul_out[881][11],mul_out[881][12],mul_out[881][13],conv_out[293]);



mul_8x8bit m2646 (image[316],filter[0],mul_out[882][11]);
mul_8x8bit m2647 (image[317],filter[1],mul_out[882][12]);
mul_8x8bit m2648 (image[318],filter[2],mul_out[882][13]);
mul_8x8bit m2649 (image[344],filter[3],mul_out[883][11]);
mul_8x8bit m2650 (image[345],filter[4],mul_out[883][12]);
mul_8x8bit m2651 (image[346],filter[5],mul_out[883][13]);
mul_8x8bit m2652 (image[372],filter[6],mul_out[884][11]);
mul_8x8bit m2653 (image[373],filter[7],mul_out[884][12]);
mul_8x8bit m2654 (image[374],filter[8],mul_out[884][13]);

adder_8bit ad294 (mul_out[882][11],mul_out[882][12],mul_out[882][13],mul_out[883][11],mul_out[883][12],mul_out[883][13],mul_out[884][11],mul_out[884][12],mul_out[884][13],conv_out[294]);



mul_8x8bit m2655 (image[317],filter[0],mul_out[885][11]);
mul_8x8bit m2656 (image[318],filter[1],mul_out[885][12]);
mul_8x8bit m2657 (image[319],filter[2],mul_out[885][13]);
mul_8x8bit m2658 (image[345],filter[3],mul_out[886][11]);
mul_8x8bit m2659 (image[346],filter[4],mul_out[886][12]);
mul_8x8bit m2660 (image[347],filter[5],mul_out[886][13]);
mul_8x8bit m2661 (image[373],filter[6],mul_out[887][11]);
mul_8x8bit m2662 (image[374],filter[7],mul_out[887][12]);
mul_8x8bit m2663 (image[375],filter[8],mul_out[887][13]);

adder_8bit ad295 (mul_out[885][11],mul_out[885][12],mul_out[885][13],mul_out[886][11],mul_out[886][12],mul_out[886][13],mul_out[887][11],mul_out[887][12],mul_out[887][13],conv_out[295]);



mul_8x8bit m2664 (image[318],filter[0],mul_out[888][11]);
mul_8x8bit m2665 (image[319],filter[1],mul_out[888][12]);
mul_8x8bit m2666 (image[320],filter[2],mul_out[888][13]);
mul_8x8bit m2667 (image[346],filter[3],mul_out[889][11]);
mul_8x8bit m2668 (image[347],filter[4],mul_out[889][12]);
mul_8x8bit m2669 (image[348],filter[5],mul_out[889][13]);
mul_8x8bit m2670 (image[374],filter[6],mul_out[890][11]);
mul_8x8bit m2671 (image[375],filter[7],mul_out[890][12]);
mul_8x8bit m2672 (image[376],filter[8],mul_out[890][13]);

adder_8bit ad296 (mul_out[888][11],mul_out[888][12],mul_out[888][13],mul_out[889][11],mul_out[889][12],mul_out[889][13],mul_out[890][11],mul_out[890][12],mul_out[890][13],conv_out[296]);



mul_8x8bit m2673 (image[319],filter[0],mul_out[891][11]);
mul_8x8bit m2674 (image[320],filter[1],mul_out[891][12]);
mul_8x8bit m2675 (image[321],filter[2],mul_out[891][13]);
mul_8x8bit m2676 (image[347],filter[3],mul_out[892][11]);
mul_8x8bit m2677 (image[348],filter[4],mul_out[892][12]);
mul_8x8bit m2678 (image[349],filter[5],mul_out[892][13]);
mul_8x8bit m2679 (image[375],filter[6],mul_out[893][11]);
mul_8x8bit m2680 (image[376],filter[7],mul_out[893][12]);
mul_8x8bit m2681 (image[377],filter[8],mul_out[893][13]);

adder_8bit ad297 (mul_out[891][11],mul_out[891][12],mul_out[891][13],mul_out[892][11],mul_out[892][12],mul_out[892][13],mul_out[893][11],mul_out[893][12],mul_out[893][13],conv_out[297]);



mul_8x8bit m2682 (image[320],filter[0],mul_out[894][11]);
mul_8x8bit m2683 (image[321],filter[1],mul_out[894][12]);
mul_8x8bit m2684 (image[322],filter[2],mul_out[894][13]);
mul_8x8bit m2685 (image[348],filter[3],mul_out[895][11]);
mul_8x8bit m2686 (image[349],filter[4],mul_out[895][12]);
mul_8x8bit m2687 (image[350],filter[5],mul_out[895][13]);
mul_8x8bit m2688 (image[376],filter[6],mul_out[896][11]);
mul_8x8bit m2689 (image[377],filter[7],mul_out[896][12]);
mul_8x8bit m2690 (image[378],filter[8],mul_out[896][13]);

adder_8bit ad298 (mul_out[894][11],mul_out[894][12],mul_out[894][13],mul_out[895][11],mul_out[895][12],mul_out[895][13],mul_out[896][11],mul_out[896][12],mul_out[896][13],conv_out[298]);



mul_8x8bit m2691 (image[321],filter[0],mul_out[897][11]);
mul_8x8bit m2692 (image[322],filter[1],mul_out[897][12]);
mul_8x8bit m2693 (image[323],filter[2],mul_out[897][13]);
mul_8x8bit m2694 (image[349],filter[3],mul_out[898][11]);
mul_8x8bit m2695 (image[350],filter[4],mul_out[898][12]);
mul_8x8bit m2696 (image[351],filter[5],mul_out[898][13]);
mul_8x8bit m2697 (image[377],filter[6],mul_out[899][11]);
mul_8x8bit m2698 (image[378],filter[7],mul_out[899][12]);
mul_8x8bit m2699 (image[379],filter[8],mul_out[899][13]);

adder_8bit ad299 (mul_out[897][11],mul_out[897][12],mul_out[897][13],mul_out[898][11],mul_out[898][12],mul_out[898][13],mul_out[899][11],mul_out[899][12],mul_out[899][13],conv_out[299]);



mul_8x8bit m2700 (image[322],filter[0],mul_out[900][11]);
mul_8x8bit m2701 (image[323],filter[1],mul_out[900][12]);
mul_8x8bit m2702 (image[324],filter[2],mul_out[900][13]);
mul_8x8bit m2703 (image[350],filter[3],mul_out[901][11]);
mul_8x8bit m2704 (image[351],filter[4],mul_out[901][12]);
mul_8x8bit m2705 (image[352],filter[5],mul_out[901][13]);
mul_8x8bit m2706 (image[378],filter[6],mul_out[902][11]);
mul_8x8bit m2707 (image[379],filter[7],mul_out[902][12]);
mul_8x8bit m2708 (image[380],filter[8],mul_out[902][13]);

adder_8bit ad300 (mul_out[900][11],mul_out[900][12],mul_out[900][13],mul_out[901][11],mul_out[901][12],mul_out[901][13],mul_out[902][11],mul_out[902][12],mul_out[902][13],conv_out[300]);



mul_8x8bit m2709 (image[323],filter[0],mul_out[903][11]);
mul_8x8bit m2710 (image[324],filter[1],mul_out[903][12]);
mul_8x8bit m2711 (image[325],filter[2],mul_out[903][13]);
mul_8x8bit m2712 (image[351],filter[3],mul_out[904][11]);
mul_8x8bit m2713 (image[352],filter[4],mul_out[904][12]);
mul_8x8bit m2714 (image[353],filter[5],mul_out[904][13]);
mul_8x8bit m2715 (image[379],filter[6],mul_out[905][11]);
mul_8x8bit m2716 (image[380],filter[7],mul_out[905][12]);
mul_8x8bit m2717 (image[381],filter[8],mul_out[905][13]);

adder_8bit ad301 (mul_out[903][11],mul_out[903][12],mul_out[903][13],mul_out[904][11],mul_out[904][12],mul_out[904][13],mul_out[905][11],mul_out[905][12],mul_out[905][13],conv_out[301]);



mul_8x8bit m2718 (image[324],filter[0],mul_out[906][11]);
mul_8x8bit m2719 (image[325],filter[1],mul_out[906][12]);
mul_8x8bit m2720 (image[326],filter[2],mul_out[906][13]);
mul_8x8bit m2721 (image[352],filter[3],mul_out[907][11]);
mul_8x8bit m2722 (image[353],filter[4],mul_out[907][12]);
mul_8x8bit m2723 (image[354],filter[5],mul_out[907][13]);
mul_8x8bit m2724 (image[380],filter[6],mul_out[908][11]);
mul_8x8bit m2725 (image[381],filter[7],mul_out[908][12]);
mul_8x8bit m2726 (image[382],filter[8],mul_out[908][13]);

adder_8bit ad302 (mul_out[906][11],mul_out[906][12],mul_out[906][13],mul_out[907][11],mul_out[907][12],mul_out[907][13],mul_out[908][11],mul_out[908][12],mul_out[908][13],conv_out[302]);



mul_8x8bit m2727 (image[325],filter[0],mul_out[909][11]);
mul_8x8bit m2728 (image[326],filter[1],mul_out[909][12]);
mul_8x8bit m2729 (image[327],filter[2],mul_out[909][13]);
mul_8x8bit m2730 (image[353],filter[3],mul_out[910][11]);
mul_8x8bit m2731 (image[354],filter[4],mul_out[910][12]);
mul_8x8bit m2732 (image[355],filter[5],mul_out[910][13]);
mul_8x8bit m2733 (image[381],filter[6],mul_out[911][11]);
mul_8x8bit m2734 (image[382],filter[7],mul_out[911][12]);
mul_8x8bit m2735 (image[383],filter[8],mul_out[911][13]);

adder_8bit ad303 (mul_out[909][11],mul_out[909][12],mul_out[909][13],mul_out[910][11],mul_out[910][12],mul_out[910][13],mul_out[911][11],mul_out[911][12],mul_out[911][13],conv_out[303]);



mul_8x8bit m2736 (image[326],filter[0],mul_out[912][11]);
mul_8x8bit m2737 (image[327],filter[1],mul_out[912][12]);
mul_8x8bit m2738 (image[328],filter[2],mul_out[912][13]);
mul_8x8bit m2739 (image[354],filter[3],mul_out[913][11]);
mul_8x8bit m2740 (image[355],filter[4],mul_out[913][12]);
mul_8x8bit m2741 (image[356],filter[5],mul_out[913][13]);
mul_8x8bit m2742 (image[382],filter[6],mul_out[914][11]);
mul_8x8bit m2743 (image[383],filter[7],mul_out[914][12]);
mul_8x8bit m2744 (image[384],filter[8],mul_out[914][13]);

adder_8bit ad304 (mul_out[912][11],mul_out[912][12],mul_out[912][13],mul_out[913][11],mul_out[913][12],mul_out[913][13],mul_out[914][11],mul_out[914][12],mul_out[914][13],conv_out[304]);



mul_8x8bit m2745 (image[327],filter[0],mul_out[915][11]);
mul_8x8bit m2746 (image[328],filter[1],mul_out[915][12]);
mul_8x8bit m2747 (image[329],filter[2],mul_out[915][13]);
mul_8x8bit m2748 (image[355],filter[3],mul_out[916][11]);
mul_8x8bit m2749 (image[356],filter[4],mul_out[916][12]);
mul_8x8bit m2750 (image[357],filter[5],mul_out[916][13]);
mul_8x8bit m2751 (image[383],filter[6],mul_out[917][11]);
mul_8x8bit m2752 (image[384],filter[7],mul_out[917][12]);
mul_8x8bit m2753 (image[385],filter[8],mul_out[917][13]);

adder_8bit ad305 (mul_out[915][11],mul_out[915][12],mul_out[915][13],mul_out[916][11],mul_out[916][12],mul_out[916][13],mul_out[917][11],mul_out[917][12],mul_out[917][13],conv_out[305]);



mul_8x8bit m2754 (image[328],filter[0],mul_out[918][11]);
mul_8x8bit m2755 (image[329],filter[1],mul_out[918][12]);
mul_8x8bit m2756 (image[330],filter[2],mul_out[918][13]);
mul_8x8bit m2757 (image[356],filter[3],mul_out[919][11]);
mul_8x8bit m2758 (image[357],filter[4],mul_out[919][12]);
mul_8x8bit m2759 (image[358],filter[5],mul_out[919][13]);
mul_8x8bit m2760 (image[384],filter[6],mul_out[920][11]);
mul_8x8bit m2761 (image[385],filter[7],mul_out[920][12]);
mul_8x8bit m2762 (image[386],filter[8],mul_out[920][13]);

adder_8bit ad306 (mul_out[918][11],mul_out[918][12],mul_out[918][13],mul_out[919][11],mul_out[919][12],mul_out[919][13],mul_out[920][11],mul_out[920][12],mul_out[920][13],conv_out[306]);



mul_8x8bit m2763 (image[329],filter[0],mul_out[921][11]);
mul_8x8bit m2764 (image[330],filter[1],mul_out[921][12]);
mul_8x8bit m2765 (image[331],filter[2],mul_out[921][13]);
mul_8x8bit m2766 (image[357],filter[3],mul_out[922][11]);
mul_8x8bit m2767 (image[358],filter[4],mul_out[922][12]);
mul_8x8bit m2768 (image[359],filter[5],mul_out[922][13]);
mul_8x8bit m2769 (image[385],filter[6],mul_out[923][11]);
mul_8x8bit m2770 (image[386],filter[7],mul_out[923][12]);
mul_8x8bit m2771 (image[387],filter[8],mul_out[923][13]);

adder_8bit ad307 (mul_out[921][11],mul_out[921][12],mul_out[921][13],mul_out[922][11],mul_out[922][12],mul_out[922][13],mul_out[923][11],mul_out[923][12],mul_out[923][13],conv_out[307]);



mul_8x8bit m2772 (image[330],filter[0],mul_out[924][11]);
mul_8x8bit m2773 (image[331],filter[1],mul_out[924][12]);
mul_8x8bit m2774 (image[332],filter[2],mul_out[924][13]);
mul_8x8bit m2775 (image[358],filter[3],mul_out[925][11]);
mul_8x8bit m2776 (image[359],filter[4],mul_out[925][12]);
mul_8x8bit m2777 (image[360],filter[5],mul_out[925][13]);
mul_8x8bit m2778 (image[386],filter[6],mul_out[926][11]);
mul_8x8bit m2779 (image[387],filter[7],mul_out[926][12]);
mul_8x8bit m2780 (image[388],filter[8],mul_out[926][13]);

adder_8bit ad308 (mul_out[924][11],mul_out[924][12],mul_out[924][13],mul_out[925][11],mul_out[925][12],mul_out[925][13],mul_out[926][11],mul_out[926][12],mul_out[926][13],conv_out[308]);



mul_8x8bit m2781 (image[331],filter[0],mul_out[927][11]);
mul_8x8bit m2782 (image[332],filter[1],mul_out[927][12]);
mul_8x8bit m2783 (image[333],filter[2],mul_out[927][13]);
mul_8x8bit m2784 (image[359],filter[3],mul_out[928][11]);
mul_8x8bit m2785 (image[360],filter[4],mul_out[928][12]);
mul_8x8bit m2786 (image[361],filter[5],mul_out[928][13]);
mul_8x8bit m2787 (image[387],filter[6],mul_out[929][11]);
mul_8x8bit m2788 (image[388],filter[7],mul_out[929][12]);
mul_8x8bit m2789 (image[389],filter[8],mul_out[929][13]);

adder_8bit ad309 (mul_out[927][11],mul_out[927][12],mul_out[927][13],mul_out[928][11],mul_out[928][12],mul_out[928][13],mul_out[929][11],mul_out[929][12],mul_out[929][13],conv_out[309]);



mul_8x8bit m2790 (image[332],filter[0],mul_out[930][11]);
mul_8x8bit m2791 (image[333],filter[1],mul_out[930][12]);
mul_8x8bit m2792 (image[334],filter[2],mul_out[930][13]);
mul_8x8bit m2793 (image[360],filter[3],mul_out[931][11]);
mul_8x8bit m2794 (image[361],filter[4],mul_out[931][12]);
mul_8x8bit m2795 (image[362],filter[5],mul_out[931][13]);
mul_8x8bit m2796 (image[388],filter[6],mul_out[932][11]);
mul_8x8bit m2797 (image[389],filter[7],mul_out[932][12]);
mul_8x8bit m2798 (image[390],filter[8],mul_out[932][13]);

adder_8bit ad310 (mul_out[930][11],mul_out[930][12],mul_out[930][13],mul_out[931][11],mul_out[931][12],mul_out[931][13],mul_out[932][11],mul_out[932][12],mul_out[932][13],conv_out[310]);



mul_8x8bit m2799 (image[333],filter[0],mul_out[933][11]);
mul_8x8bit m2800 (image[334],filter[1],mul_out[933][12]);
mul_8x8bit m2801 (image[335],filter[2],mul_out[933][13]);
mul_8x8bit m2802 (image[361],filter[3],mul_out[934][11]);
mul_8x8bit m2803 (image[362],filter[4],mul_out[934][12]);
mul_8x8bit m2804 (image[363],filter[5],mul_out[934][13]);
mul_8x8bit m2805 (image[389],filter[6],mul_out[935][11]);
mul_8x8bit m2806 (image[390],filter[7],mul_out[935][12]);
mul_8x8bit m2807 (image[391],filter[8],mul_out[935][13]);

adder_8bit ad311 (mul_out[933][11],mul_out[933][12],mul_out[933][13],mul_out[934][11],mul_out[934][12],mul_out[934][13],mul_out[935][11],mul_out[935][12],mul_out[935][13],conv_out[311]);



mul_8x8bit m2808 (image[336],filter[0],mul_out[936][12]);
mul_8x8bit m2809 (image[337],filter[1],mul_out[936][13]);
mul_8x8bit m2810 (image[338],filter[2],mul_out[936][14]);
mul_8x8bit m2811 (image[364],filter[3],mul_out[937][12]);
mul_8x8bit m2812 (image[365],filter[4],mul_out[937][13]);
mul_8x8bit m2813 (image[366],filter[5],mul_out[937][14]);
mul_8x8bit m2814 (image[392],filter[6],mul_out[938][12]);
mul_8x8bit m2815 (image[393],filter[7],mul_out[938][13]);
mul_8x8bit m2816 (image[394],filter[8],mul_out[938][14]);

adder_8bit ad312 (mul_out[936][12],mul_out[936][13],mul_out[936][14],mul_out[937][12],mul_out[937][13],mul_out[937][14],mul_out[938][12],mul_out[938][13],mul_out[938][14],conv_out[312]);



mul_8x8bit m2817 (image[337],filter[0],mul_out[939][12]);
mul_8x8bit m2818 (image[338],filter[1],mul_out[939][13]);
mul_8x8bit m2819 (image[339],filter[2],mul_out[939][14]);
mul_8x8bit m2820 (image[365],filter[3],mul_out[940][12]);
mul_8x8bit m2821 (image[366],filter[4],mul_out[940][13]);
mul_8x8bit m2822 (image[367],filter[5],mul_out[940][14]);
mul_8x8bit m2823 (image[393],filter[6],mul_out[941][12]);
mul_8x8bit m2824 (image[394],filter[7],mul_out[941][13]);
mul_8x8bit m2825 (image[395],filter[8],mul_out[941][14]);

adder_8bit ad313 (mul_out[939][12],mul_out[939][13],mul_out[939][14],mul_out[940][12],mul_out[940][13],mul_out[940][14],mul_out[941][12],mul_out[941][13],mul_out[941][14],conv_out[313]);



mul_8x8bit m2826 (image[338],filter[0],mul_out[942][12]);
mul_8x8bit m2827 (image[339],filter[1],mul_out[942][13]);
mul_8x8bit m2828 (image[340],filter[2],mul_out[942][14]);
mul_8x8bit m2829 (image[366],filter[3],mul_out[943][12]);
mul_8x8bit m2830 (image[367],filter[4],mul_out[943][13]);
mul_8x8bit m2831 (image[368],filter[5],mul_out[943][14]);
mul_8x8bit m2832 (image[394],filter[6],mul_out[944][12]);
mul_8x8bit m2833 (image[395],filter[7],mul_out[944][13]);
mul_8x8bit m2834 (image[396],filter[8],mul_out[944][14]);

adder_8bit ad314 (mul_out[942][12],mul_out[942][13],mul_out[942][14],mul_out[943][12],mul_out[943][13],mul_out[943][14],mul_out[944][12],mul_out[944][13],mul_out[944][14],conv_out[314]);



mul_8x8bit m2835 (image[339],filter[0],mul_out[945][12]);
mul_8x8bit m2836 (image[340],filter[1],mul_out[945][13]);
mul_8x8bit m2837 (image[341],filter[2],mul_out[945][14]);
mul_8x8bit m2838 (image[367],filter[3],mul_out[946][12]);
mul_8x8bit m2839 (image[368],filter[4],mul_out[946][13]);
mul_8x8bit m2840 (image[369],filter[5],mul_out[946][14]);
mul_8x8bit m2841 (image[395],filter[6],mul_out[947][12]);
mul_8x8bit m2842 (image[396],filter[7],mul_out[947][13]);
mul_8x8bit m2843 (image[397],filter[8],mul_out[947][14]);

adder_8bit ad315 (mul_out[945][12],mul_out[945][13],mul_out[945][14],mul_out[946][12],mul_out[946][13],mul_out[946][14],mul_out[947][12],mul_out[947][13],mul_out[947][14],conv_out[315]);



mul_8x8bit m2844 (image[340],filter[0],mul_out[948][12]);
mul_8x8bit m2845 (image[341],filter[1],mul_out[948][13]);
mul_8x8bit m2846 (image[342],filter[2],mul_out[948][14]);
mul_8x8bit m2847 (image[368],filter[3],mul_out[949][12]);
mul_8x8bit m2848 (image[369],filter[4],mul_out[949][13]);
mul_8x8bit m2849 (image[370],filter[5],mul_out[949][14]);
mul_8x8bit m2850 (image[396],filter[6],mul_out[950][12]);
mul_8x8bit m2851 (image[397],filter[7],mul_out[950][13]);
mul_8x8bit m2852 (image[398],filter[8],mul_out[950][14]);

adder_8bit ad316 (mul_out[948][12],mul_out[948][13],mul_out[948][14],mul_out[949][12],mul_out[949][13],mul_out[949][14],mul_out[950][12],mul_out[950][13],mul_out[950][14],conv_out[316]);



mul_8x8bit m2853 (image[341],filter[0],mul_out[951][12]);
mul_8x8bit m2854 (image[342],filter[1],mul_out[951][13]);
mul_8x8bit m2855 (image[343],filter[2],mul_out[951][14]);
mul_8x8bit m2856 (image[369],filter[3],mul_out[952][12]);
mul_8x8bit m2857 (image[370],filter[4],mul_out[952][13]);
mul_8x8bit m2858 (image[371],filter[5],mul_out[952][14]);
mul_8x8bit m2859 (image[397],filter[6],mul_out[953][12]);
mul_8x8bit m2860 (image[398],filter[7],mul_out[953][13]);
mul_8x8bit m2861 (image[399],filter[8],mul_out[953][14]);

adder_8bit ad317 (mul_out[951][12],mul_out[951][13],mul_out[951][14],mul_out[952][12],mul_out[952][13],mul_out[952][14],mul_out[953][12],mul_out[953][13],mul_out[953][14],conv_out[317]);



mul_8x8bit m2862 (image[342],filter[0],mul_out[954][12]);
mul_8x8bit m2863 (image[343],filter[1],mul_out[954][13]);
mul_8x8bit m2864 (image[344],filter[2],mul_out[954][14]);
mul_8x8bit m2865 (image[370],filter[3],mul_out[955][12]);
mul_8x8bit m2866 (image[371],filter[4],mul_out[955][13]);
mul_8x8bit m2867 (image[372],filter[5],mul_out[955][14]);
mul_8x8bit m2868 (image[398],filter[6],mul_out[956][12]);
mul_8x8bit m2869 (image[399],filter[7],mul_out[956][13]);
mul_8x8bit m2870 (image[400],filter[8],mul_out[956][14]);

adder_8bit ad318 (mul_out[954][12],mul_out[954][13],mul_out[954][14],mul_out[955][12],mul_out[955][13],mul_out[955][14],mul_out[956][12],mul_out[956][13],mul_out[956][14],conv_out[318]);



mul_8x8bit m2871 (image[343],filter[0],mul_out[957][12]);
mul_8x8bit m2872 (image[344],filter[1],mul_out[957][13]);
mul_8x8bit m2873 (image[345],filter[2],mul_out[957][14]);
mul_8x8bit m2874 (image[371],filter[3],mul_out[958][12]);
mul_8x8bit m2875 (image[372],filter[4],mul_out[958][13]);
mul_8x8bit m2876 (image[373],filter[5],mul_out[958][14]);
mul_8x8bit m2877 (image[399],filter[6],mul_out[959][12]);
mul_8x8bit m2878 (image[400],filter[7],mul_out[959][13]);
mul_8x8bit m2879 (image[401],filter[8],mul_out[959][14]);

adder_8bit ad319 (mul_out[957][12],mul_out[957][13],mul_out[957][14],mul_out[958][12],mul_out[958][13],mul_out[958][14],mul_out[959][12],mul_out[959][13],mul_out[959][14],conv_out[319]);



mul_8x8bit m2880 (image[344],filter[0],mul_out[960][12]);
mul_8x8bit m2881 (image[345],filter[1],mul_out[960][13]);
mul_8x8bit m2882 (image[346],filter[2],mul_out[960][14]);
mul_8x8bit m2883 (image[372],filter[3],mul_out[961][12]);
mul_8x8bit m2884 (image[373],filter[4],mul_out[961][13]);
mul_8x8bit m2885 (image[374],filter[5],mul_out[961][14]);
mul_8x8bit m2886 (image[400],filter[6],mul_out[962][12]);
mul_8x8bit m2887 (image[401],filter[7],mul_out[962][13]);
mul_8x8bit m2888 (image[402],filter[8],mul_out[962][14]);

adder_8bit ad320 (mul_out[960][12],mul_out[960][13],mul_out[960][14],mul_out[961][12],mul_out[961][13],mul_out[961][14],mul_out[962][12],mul_out[962][13],mul_out[962][14],conv_out[320]);



mul_8x8bit m2889 (image[345],filter[0],mul_out[963][12]);
mul_8x8bit m2890 (image[346],filter[1],mul_out[963][13]);
mul_8x8bit m2891 (image[347],filter[2],mul_out[963][14]);
mul_8x8bit m2892 (image[373],filter[3],mul_out[964][12]);
mul_8x8bit m2893 (image[374],filter[4],mul_out[964][13]);
mul_8x8bit m2894 (image[375],filter[5],mul_out[964][14]);
mul_8x8bit m2895 (image[401],filter[6],mul_out[965][12]);
mul_8x8bit m2896 (image[402],filter[7],mul_out[965][13]);
mul_8x8bit m2897 (image[403],filter[8],mul_out[965][14]);

adder_8bit ad321 (mul_out[963][12],mul_out[963][13],mul_out[963][14],mul_out[964][12],mul_out[964][13],mul_out[964][14],mul_out[965][12],mul_out[965][13],mul_out[965][14],conv_out[321]);



mul_8x8bit m2898 (image[346],filter[0],mul_out[966][12]);
mul_8x8bit m2899 (image[347],filter[1],mul_out[966][13]);
mul_8x8bit m2900 (image[348],filter[2],mul_out[966][14]);
mul_8x8bit m2901 (image[374],filter[3],mul_out[967][12]);
mul_8x8bit m2902 (image[375],filter[4],mul_out[967][13]);
mul_8x8bit m2903 (image[376],filter[5],mul_out[967][14]);
mul_8x8bit m2904 (image[402],filter[6],mul_out[968][12]);
mul_8x8bit m2905 (image[403],filter[7],mul_out[968][13]);
mul_8x8bit m2906 (image[404],filter[8],mul_out[968][14]);

adder_8bit ad322 (mul_out[966][12],mul_out[966][13],mul_out[966][14],mul_out[967][12],mul_out[967][13],mul_out[967][14],mul_out[968][12],mul_out[968][13],mul_out[968][14],conv_out[322]);



mul_8x8bit m2907 (image[347],filter[0],mul_out[969][12]);
mul_8x8bit m2908 (image[348],filter[1],mul_out[969][13]);
mul_8x8bit m2909 (image[349],filter[2],mul_out[969][14]);
mul_8x8bit m2910 (image[375],filter[3],mul_out[970][12]);
mul_8x8bit m2911 (image[376],filter[4],mul_out[970][13]);
mul_8x8bit m2912 (image[377],filter[5],mul_out[970][14]);
mul_8x8bit m2913 (image[403],filter[6],mul_out[971][12]);
mul_8x8bit m2914 (image[404],filter[7],mul_out[971][13]);
mul_8x8bit m2915 (image[405],filter[8],mul_out[971][14]);

adder_8bit ad323 (mul_out[969][12],mul_out[969][13],mul_out[969][14],mul_out[970][12],mul_out[970][13],mul_out[970][14],mul_out[971][12],mul_out[971][13],mul_out[971][14],conv_out[323]);



mul_8x8bit m2916 (image[348],filter[0],mul_out[972][12]);
mul_8x8bit m2917 (image[349],filter[1],mul_out[972][13]);
mul_8x8bit m2918 (image[350],filter[2],mul_out[972][14]);
mul_8x8bit m2919 (image[376],filter[3],mul_out[973][12]);
mul_8x8bit m2920 (image[377],filter[4],mul_out[973][13]);
mul_8x8bit m2921 (image[378],filter[5],mul_out[973][14]);
mul_8x8bit m2922 (image[404],filter[6],mul_out[974][12]);
mul_8x8bit m2923 (image[405],filter[7],mul_out[974][13]);
mul_8x8bit m2924 (image[406],filter[8],mul_out[974][14]);

adder_8bit ad324 (mul_out[972][12],mul_out[972][13],mul_out[972][14],mul_out[973][12],mul_out[973][13],mul_out[973][14],mul_out[974][12],mul_out[974][13],mul_out[974][14],conv_out[324]);



mul_8x8bit m2925 (image[349],filter[0],mul_out[975][12]);
mul_8x8bit m2926 (image[350],filter[1],mul_out[975][13]);
mul_8x8bit m2927 (image[351],filter[2],mul_out[975][14]);
mul_8x8bit m2928 (image[377],filter[3],mul_out[976][12]);
mul_8x8bit m2929 (image[378],filter[4],mul_out[976][13]);
mul_8x8bit m2930 (image[379],filter[5],mul_out[976][14]);
mul_8x8bit m2931 (image[405],filter[6],mul_out[977][12]);
mul_8x8bit m2932 (image[406],filter[7],mul_out[977][13]);
mul_8x8bit m2933 (image[407],filter[8],mul_out[977][14]);

adder_8bit ad325 (mul_out[975][12],mul_out[975][13],mul_out[975][14],mul_out[976][12],mul_out[976][13],mul_out[976][14],mul_out[977][12],mul_out[977][13],mul_out[977][14],conv_out[325]);



mul_8x8bit m2934 (image[350],filter[0],mul_out[978][12]);
mul_8x8bit m2935 (image[351],filter[1],mul_out[978][13]);
mul_8x8bit m2936 (image[352],filter[2],mul_out[978][14]);
mul_8x8bit m2937 (image[378],filter[3],mul_out[979][12]);
mul_8x8bit m2938 (image[379],filter[4],mul_out[979][13]);
mul_8x8bit m2939 (image[380],filter[5],mul_out[979][14]);
mul_8x8bit m2940 (image[406],filter[6],mul_out[980][12]);
mul_8x8bit m2941 (image[407],filter[7],mul_out[980][13]);
mul_8x8bit m2942 (image[408],filter[8],mul_out[980][14]);

adder_8bit ad326 (mul_out[978][12],mul_out[978][13],mul_out[978][14],mul_out[979][12],mul_out[979][13],mul_out[979][14],mul_out[980][12],mul_out[980][13],mul_out[980][14],conv_out[326]);



mul_8x8bit m2943 (image[351],filter[0],mul_out[981][12]);
mul_8x8bit m2944 (image[352],filter[1],mul_out[981][13]);
mul_8x8bit m2945 (image[353],filter[2],mul_out[981][14]);
mul_8x8bit m2946 (image[379],filter[3],mul_out[982][12]);
mul_8x8bit m2947 (image[380],filter[4],mul_out[982][13]);
mul_8x8bit m2948 (image[381],filter[5],mul_out[982][14]);
mul_8x8bit m2949 (image[407],filter[6],mul_out[983][12]);
mul_8x8bit m2950 (image[408],filter[7],mul_out[983][13]);
mul_8x8bit m2951 (image[409],filter[8],mul_out[983][14]);

adder_8bit ad327 (mul_out[981][12],mul_out[981][13],mul_out[981][14],mul_out[982][12],mul_out[982][13],mul_out[982][14],mul_out[983][12],mul_out[983][13],mul_out[983][14],conv_out[327]);



mul_8x8bit m2952 (image[352],filter[0],mul_out[984][12]);
mul_8x8bit m2953 (image[353],filter[1],mul_out[984][13]);
mul_8x8bit m2954 (image[354],filter[2],mul_out[984][14]);
mul_8x8bit m2955 (image[380],filter[3],mul_out[985][12]);
mul_8x8bit m2956 (image[381],filter[4],mul_out[985][13]);
mul_8x8bit m2957 (image[382],filter[5],mul_out[985][14]);
mul_8x8bit m2958 (image[408],filter[6],mul_out[986][12]);
mul_8x8bit m2959 (image[409],filter[7],mul_out[986][13]);
mul_8x8bit m2960 (image[410],filter[8],mul_out[986][14]);

adder_8bit ad328 (mul_out[984][12],mul_out[984][13],mul_out[984][14],mul_out[985][12],mul_out[985][13],mul_out[985][14],mul_out[986][12],mul_out[986][13],mul_out[986][14],conv_out[328]);



mul_8x8bit m2961 (image[353],filter[0],mul_out[987][12]);
mul_8x8bit m2962 (image[354],filter[1],mul_out[987][13]);
mul_8x8bit m2963 (image[355],filter[2],mul_out[987][14]);
mul_8x8bit m2964 (image[381],filter[3],mul_out[988][12]);
mul_8x8bit m2965 (image[382],filter[4],mul_out[988][13]);
mul_8x8bit m2966 (image[383],filter[5],mul_out[988][14]);
mul_8x8bit m2967 (image[409],filter[6],mul_out[989][12]);
mul_8x8bit m2968 (image[410],filter[7],mul_out[989][13]);
mul_8x8bit m2969 (image[411],filter[8],mul_out[989][14]);

adder_8bit ad329 (mul_out[987][12],mul_out[987][13],mul_out[987][14],mul_out[988][12],mul_out[988][13],mul_out[988][14],mul_out[989][12],mul_out[989][13],mul_out[989][14],conv_out[329]);



mul_8x8bit m2970 (image[354],filter[0],mul_out[990][12]);
mul_8x8bit m2971 (image[355],filter[1],mul_out[990][13]);
mul_8x8bit m2972 (image[356],filter[2],mul_out[990][14]);
mul_8x8bit m2973 (image[382],filter[3],mul_out[991][12]);
mul_8x8bit m2974 (image[383],filter[4],mul_out[991][13]);
mul_8x8bit m2975 (image[384],filter[5],mul_out[991][14]);
mul_8x8bit m2976 (image[410],filter[6],mul_out[992][12]);
mul_8x8bit m2977 (image[411],filter[7],mul_out[992][13]);
mul_8x8bit m2978 (image[412],filter[8],mul_out[992][14]);

adder_8bit ad330 (mul_out[990][12],mul_out[990][13],mul_out[990][14],mul_out[991][12],mul_out[991][13],mul_out[991][14],mul_out[992][12],mul_out[992][13],mul_out[992][14],conv_out[330]);



mul_8x8bit m2979 (image[355],filter[0],mul_out[993][12]);
mul_8x8bit m2980 (image[356],filter[1],mul_out[993][13]);
mul_8x8bit m2981 (image[357],filter[2],mul_out[993][14]);
mul_8x8bit m2982 (image[383],filter[3],mul_out[994][12]);
mul_8x8bit m2983 (image[384],filter[4],mul_out[994][13]);
mul_8x8bit m2984 (image[385],filter[5],mul_out[994][14]);
mul_8x8bit m2985 (image[411],filter[6],mul_out[995][12]);
mul_8x8bit m2986 (image[412],filter[7],mul_out[995][13]);
mul_8x8bit m2987 (image[413],filter[8],mul_out[995][14]);

adder_8bit ad331 (mul_out[993][12],mul_out[993][13],mul_out[993][14],mul_out[994][12],mul_out[994][13],mul_out[994][14],mul_out[995][12],mul_out[995][13],mul_out[995][14],conv_out[331]);



mul_8x8bit m2988 (image[356],filter[0],mul_out[996][12]);
mul_8x8bit m2989 (image[357],filter[1],mul_out[996][13]);
mul_8x8bit m2990 (image[358],filter[2],mul_out[996][14]);
mul_8x8bit m2991 (image[384],filter[3],mul_out[997][12]);
mul_8x8bit m2992 (image[385],filter[4],mul_out[997][13]);
mul_8x8bit m2993 (image[386],filter[5],mul_out[997][14]);
mul_8x8bit m2994 (image[412],filter[6],mul_out[998][12]);
mul_8x8bit m2995 (image[413],filter[7],mul_out[998][13]);
mul_8x8bit m2996 (image[414],filter[8],mul_out[998][14]);

adder_8bit ad332 (mul_out[996][12],mul_out[996][13],mul_out[996][14],mul_out[997][12],mul_out[997][13],mul_out[997][14],mul_out[998][12],mul_out[998][13],mul_out[998][14],conv_out[332]);



mul_8x8bit m2997 (image[357],filter[0],mul_out[999][12]);
mul_8x8bit m2998 (image[358],filter[1],mul_out[999][13]);
mul_8x8bit m2999 (image[359],filter[2],mul_out[999][14]);
mul_8x8bit m3000 (image[385],filter[3],mul_out[1000][12]);
mul_8x8bit m3001 (image[386],filter[4],mul_out[1000][13]);
mul_8x8bit m3002 (image[387],filter[5],mul_out[1000][14]);
mul_8x8bit m3003 (image[413],filter[6],mul_out[1001][12]);
mul_8x8bit m3004 (image[414],filter[7],mul_out[1001][13]);
mul_8x8bit m3005 (image[415],filter[8],mul_out[1001][14]);

adder_8bit ad333 (mul_out[999][12],mul_out[999][13],mul_out[999][14],mul_out[1000][12],mul_out[1000][13],mul_out[1000][14],mul_out[1001][12],mul_out[1001][13],mul_out[1001][14],conv_out[333]);



mul_8x8bit m3006 (image[358],filter[0],mul_out[1002][12]);
mul_8x8bit m3007 (image[359],filter[1],mul_out[1002][13]);
mul_8x8bit m3008 (image[360],filter[2],mul_out[1002][14]);
mul_8x8bit m3009 (image[386],filter[3],mul_out[1003][12]);
mul_8x8bit m3010 (image[387],filter[4],mul_out[1003][13]);
mul_8x8bit m3011 (image[388],filter[5],mul_out[1003][14]);
mul_8x8bit m3012 (image[414],filter[6],mul_out[1004][12]);
mul_8x8bit m3013 (image[415],filter[7],mul_out[1004][13]);
mul_8x8bit m3014 (image[416],filter[8],mul_out[1004][14]);

adder_8bit ad334 (mul_out[1002][12],mul_out[1002][13],mul_out[1002][14],mul_out[1003][12],mul_out[1003][13],mul_out[1003][14],mul_out[1004][12],mul_out[1004][13],mul_out[1004][14],conv_out[334]);



mul_8x8bit m3015 (image[359],filter[0],mul_out[1005][12]);
mul_8x8bit m3016 (image[360],filter[1],mul_out[1005][13]);
mul_8x8bit m3017 (image[361],filter[2],mul_out[1005][14]);
mul_8x8bit m3018 (image[387],filter[3],mul_out[1006][12]);
mul_8x8bit m3019 (image[388],filter[4],mul_out[1006][13]);
mul_8x8bit m3020 (image[389],filter[5],mul_out[1006][14]);
mul_8x8bit m3021 (image[415],filter[6],mul_out[1007][12]);
mul_8x8bit m3022 (image[416],filter[7],mul_out[1007][13]);
mul_8x8bit m3023 (image[417],filter[8],mul_out[1007][14]);

adder_8bit ad335 (mul_out[1005][12],mul_out[1005][13],mul_out[1005][14],mul_out[1006][12],mul_out[1006][13],mul_out[1006][14],mul_out[1007][12],mul_out[1007][13],mul_out[1007][14],conv_out[335]);



mul_8x8bit m3024 (image[360],filter[0],mul_out[1008][12]);
mul_8x8bit m3025 (image[361],filter[1],mul_out[1008][13]);
mul_8x8bit m3026 (image[362],filter[2],mul_out[1008][14]);
mul_8x8bit m3027 (image[388],filter[3],mul_out[1009][12]);
mul_8x8bit m3028 (image[389],filter[4],mul_out[1009][13]);
mul_8x8bit m3029 (image[390],filter[5],mul_out[1009][14]);
mul_8x8bit m3030 (image[416],filter[6],mul_out[1010][12]);
mul_8x8bit m3031 (image[417],filter[7],mul_out[1010][13]);
mul_8x8bit m3032 (image[418],filter[8],mul_out[1010][14]);

adder_8bit ad336 (mul_out[1008][12],mul_out[1008][13],mul_out[1008][14],mul_out[1009][12],mul_out[1009][13],mul_out[1009][14],mul_out[1010][12],mul_out[1010][13],mul_out[1010][14],conv_out[336]);



mul_8x8bit m3033 (image[361],filter[0],mul_out[1011][12]);
mul_8x8bit m3034 (image[362],filter[1],mul_out[1011][13]);
mul_8x8bit m3035 (image[363],filter[2],mul_out[1011][14]);
mul_8x8bit m3036 (image[389],filter[3],mul_out[1012][12]);
mul_8x8bit m3037 (image[390],filter[4],mul_out[1012][13]);
mul_8x8bit m3038 (image[391],filter[5],mul_out[1012][14]);
mul_8x8bit m3039 (image[417],filter[6],mul_out[1013][12]);
mul_8x8bit m3040 (image[418],filter[7],mul_out[1013][13]);
mul_8x8bit m3041 (image[419],filter[8],mul_out[1013][14]);

adder_8bit ad337 (mul_out[1011][12],mul_out[1011][13],mul_out[1011][14],mul_out[1012][12],mul_out[1012][13],mul_out[1012][14],mul_out[1013][12],mul_out[1013][13],mul_out[1013][14],conv_out[337]);



mul_8x8bit m3042 (image[364],filter[0],mul_out[1014][13]);
mul_8x8bit m3043 (image[365],filter[1],mul_out[1014][14]);
mul_8x8bit m3044 (image[366],filter[2],mul_out[1014][15]);
mul_8x8bit m3045 (image[392],filter[3],mul_out[1015][13]);
mul_8x8bit m3046 (image[393],filter[4],mul_out[1015][14]);
mul_8x8bit m3047 (image[394],filter[5],mul_out[1015][15]);
mul_8x8bit m3048 (image[420],filter[6],mul_out[1016][13]);
mul_8x8bit m3049 (image[421],filter[7],mul_out[1016][14]);
mul_8x8bit m3050 (image[422],filter[8],mul_out[1016][15]);

adder_8bit ad338 (mul_out[1014][13],mul_out[1014][14],mul_out[1014][15],mul_out[1015][13],mul_out[1015][14],mul_out[1015][15],mul_out[1016][13],mul_out[1016][14],mul_out[1016][15],conv_out[338]);



mul_8x8bit m3051 (image[365],filter[0],mul_out[1017][13]);
mul_8x8bit m3052 (image[366],filter[1],mul_out[1017][14]);
mul_8x8bit m3053 (image[367],filter[2],mul_out[1017][15]);
mul_8x8bit m3054 (image[393],filter[3],mul_out[1018][13]);
mul_8x8bit m3055 (image[394],filter[4],mul_out[1018][14]);
mul_8x8bit m3056 (image[395],filter[5],mul_out[1018][15]);
mul_8x8bit m3057 (image[421],filter[6],mul_out[1019][13]);
mul_8x8bit m3058 (image[422],filter[7],mul_out[1019][14]);
mul_8x8bit m3059 (image[423],filter[8],mul_out[1019][15]);

adder_8bit ad339 (mul_out[1017][13],mul_out[1017][14],mul_out[1017][15],mul_out[1018][13],mul_out[1018][14],mul_out[1018][15],mul_out[1019][13],mul_out[1019][14],mul_out[1019][15],conv_out[339]);



mul_8x8bit m3060 (image[366],filter[0],mul_out[1020][13]);
mul_8x8bit m3061 (image[367],filter[1],mul_out[1020][14]);
mul_8x8bit m3062 (image[368],filter[2],mul_out[1020][15]);
mul_8x8bit m3063 (image[394],filter[3],mul_out[1021][13]);
mul_8x8bit m3064 (image[395],filter[4],mul_out[1021][14]);
mul_8x8bit m3065 (image[396],filter[5],mul_out[1021][15]);
mul_8x8bit m3066 (image[422],filter[6],mul_out[1022][13]);
mul_8x8bit m3067 (image[423],filter[7],mul_out[1022][14]);
mul_8x8bit m3068 (image[424],filter[8],mul_out[1022][15]);

adder_8bit ad340 (mul_out[1020][13],mul_out[1020][14],mul_out[1020][15],mul_out[1021][13],mul_out[1021][14],mul_out[1021][15],mul_out[1022][13],mul_out[1022][14],mul_out[1022][15],conv_out[340]);



mul_8x8bit m3069 (image[367],filter[0],mul_out[1023][13]);
mul_8x8bit m3070 (image[368],filter[1],mul_out[1023][14]);
mul_8x8bit m3071 (image[369],filter[2],mul_out[1023][15]);
mul_8x8bit m3072 (image[395],filter[3],mul_out[1024][13]);
mul_8x8bit m3073 (image[396],filter[4],mul_out[1024][14]);
mul_8x8bit m3074 (image[397],filter[5],mul_out[1024][15]);
mul_8x8bit m3075 (image[423],filter[6],mul_out[1025][13]);
mul_8x8bit m3076 (image[424],filter[7],mul_out[1025][14]);
mul_8x8bit m3077 (image[425],filter[8],mul_out[1025][15]);

adder_8bit ad341 (mul_out[1023][13],mul_out[1023][14],mul_out[1023][15],mul_out[1024][13],mul_out[1024][14],mul_out[1024][15],mul_out[1025][13],mul_out[1025][14],mul_out[1025][15],conv_out[341]);



mul_8x8bit m3078 (image[368],filter[0],mul_out[1026][13]);
mul_8x8bit m3079 (image[369],filter[1],mul_out[1026][14]);
mul_8x8bit m3080 (image[370],filter[2],mul_out[1026][15]);
mul_8x8bit m3081 (image[396],filter[3],mul_out[1027][13]);
mul_8x8bit m3082 (image[397],filter[4],mul_out[1027][14]);
mul_8x8bit m3083 (image[398],filter[5],mul_out[1027][15]);
mul_8x8bit m3084 (image[424],filter[6],mul_out[1028][13]);
mul_8x8bit m3085 (image[425],filter[7],mul_out[1028][14]);
mul_8x8bit m3086 (image[426],filter[8],mul_out[1028][15]);

adder_8bit ad342 (mul_out[1026][13],mul_out[1026][14],mul_out[1026][15],mul_out[1027][13],mul_out[1027][14],mul_out[1027][15],mul_out[1028][13],mul_out[1028][14],mul_out[1028][15],conv_out[342]);



mul_8x8bit m3087 (image[369],filter[0],mul_out[1029][13]);
mul_8x8bit m3088 (image[370],filter[1],mul_out[1029][14]);
mul_8x8bit m3089 (image[371],filter[2],mul_out[1029][15]);
mul_8x8bit m3090 (image[397],filter[3],mul_out[1030][13]);
mul_8x8bit m3091 (image[398],filter[4],mul_out[1030][14]);
mul_8x8bit m3092 (image[399],filter[5],mul_out[1030][15]);
mul_8x8bit m3093 (image[425],filter[6],mul_out[1031][13]);
mul_8x8bit m3094 (image[426],filter[7],mul_out[1031][14]);
mul_8x8bit m3095 (image[427],filter[8],mul_out[1031][15]);

adder_8bit ad343 (mul_out[1029][13],mul_out[1029][14],mul_out[1029][15],mul_out[1030][13],mul_out[1030][14],mul_out[1030][15],mul_out[1031][13],mul_out[1031][14],mul_out[1031][15],conv_out[343]);



mul_8x8bit m3096 (image[370],filter[0],mul_out[1032][13]);
mul_8x8bit m3097 (image[371],filter[1],mul_out[1032][14]);
mul_8x8bit m3098 (image[372],filter[2],mul_out[1032][15]);
mul_8x8bit m3099 (image[398],filter[3],mul_out[1033][13]);
mul_8x8bit m3100 (image[399],filter[4],mul_out[1033][14]);
mul_8x8bit m3101 (image[400],filter[5],mul_out[1033][15]);
mul_8x8bit m3102 (image[426],filter[6],mul_out[1034][13]);
mul_8x8bit m3103 (image[427],filter[7],mul_out[1034][14]);
mul_8x8bit m3104 (image[428],filter[8],mul_out[1034][15]);

adder_8bit ad344 (mul_out[1032][13],mul_out[1032][14],mul_out[1032][15],mul_out[1033][13],mul_out[1033][14],mul_out[1033][15],mul_out[1034][13],mul_out[1034][14],mul_out[1034][15],conv_out[344]);



mul_8x8bit m3105 (image[371],filter[0],mul_out[1035][13]);
mul_8x8bit m3106 (image[372],filter[1],mul_out[1035][14]);
mul_8x8bit m3107 (image[373],filter[2],mul_out[1035][15]);
mul_8x8bit m3108 (image[399],filter[3],mul_out[1036][13]);
mul_8x8bit m3109 (image[400],filter[4],mul_out[1036][14]);
mul_8x8bit m3110 (image[401],filter[5],mul_out[1036][15]);
mul_8x8bit m3111 (image[427],filter[6],mul_out[1037][13]);
mul_8x8bit m3112 (image[428],filter[7],mul_out[1037][14]);
mul_8x8bit m3113 (image[429],filter[8],mul_out[1037][15]);

adder_8bit ad345 (mul_out[1035][13],mul_out[1035][14],mul_out[1035][15],mul_out[1036][13],mul_out[1036][14],mul_out[1036][15],mul_out[1037][13],mul_out[1037][14],mul_out[1037][15],conv_out[345]);



mul_8x8bit m3114 (image[372],filter[0],mul_out[1038][13]);
mul_8x8bit m3115 (image[373],filter[1],mul_out[1038][14]);
mul_8x8bit m3116 (image[374],filter[2],mul_out[1038][15]);
mul_8x8bit m3117 (image[400],filter[3],mul_out[1039][13]);
mul_8x8bit m3118 (image[401],filter[4],mul_out[1039][14]);
mul_8x8bit m3119 (image[402],filter[5],mul_out[1039][15]);
mul_8x8bit m3120 (image[428],filter[6],mul_out[1040][13]);
mul_8x8bit m3121 (image[429],filter[7],mul_out[1040][14]);
mul_8x8bit m3122 (image[430],filter[8],mul_out[1040][15]);

adder_8bit ad346 (mul_out[1038][13],mul_out[1038][14],mul_out[1038][15],mul_out[1039][13],mul_out[1039][14],mul_out[1039][15],mul_out[1040][13],mul_out[1040][14],mul_out[1040][15],conv_out[346]);



mul_8x8bit m3123 (image[373],filter[0],mul_out[1041][13]);
mul_8x8bit m3124 (image[374],filter[1],mul_out[1041][14]);
mul_8x8bit m3125 (image[375],filter[2],mul_out[1041][15]);
mul_8x8bit m3126 (image[401],filter[3],mul_out[1042][13]);
mul_8x8bit m3127 (image[402],filter[4],mul_out[1042][14]);
mul_8x8bit m3128 (image[403],filter[5],mul_out[1042][15]);
mul_8x8bit m3129 (image[429],filter[6],mul_out[1043][13]);
mul_8x8bit m3130 (image[430],filter[7],mul_out[1043][14]);
mul_8x8bit m3131 (image[431],filter[8],mul_out[1043][15]);

adder_8bit ad347 (mul_out[1041][13],mul_out[1041][14],mul_out[1041][15],mul_out[1042][13],mul_out[1042][14],mul_out[1042][15],mul_out[1043][13],mul_out[1043][14],mul_out[1043][15],conv_out[347]);



mul_8x8bit m3132 (image[374],filter[0],mul_out[1044][13]);
mul_8x8bit m3133 (image[375],filter[1],mul_out[1044][14]);
mul_8x8bit m3134 (image[376],filter[2],mul_out[1044][15]);
mul_8x8bit m3135 (image[402],filter[3],mul_out[1045][13]);
mul_8x8bit m3136 (image[403],filter[4],mul_out[1045][14]);
mul_8x8bit m3137 (image[404],filter[5],mul_out[1045][15]);
mul_8x8bit m3138 (image[430],filter[6],mul_out[1046][13]);
mul_8x8bit m3139 (image[431],filter[7],mul_out[1046][14]);
mul_8x8bit m3140 (image[432],filter[8],mul_out[1046][15]);

adder_8bit ad348 (mul_out[1044][13],mul_out[1044][14],mul_out[1044][15],mul_out[1045][13],mul_out[1045][14],mul_out[1045][15],mul_out[1046][13],mul_out[1046][14],mul_out[1046][15],conv_out[348]);



mul_8x8bit m3141 (image[375],filter[0],mul_out[1047][13]);
mul_8x8bit m3142 (image[376],filter[1],mul_out[1047][14]);
mul_8x8bit m3143 (image[377],filter[2],mul_out[1047][15]);
mul_8x8bit m3144 (image[403],filter[3],mul_out[1048][13]);
mul_8x8bit m3145 (image[404],filter[4],mul_out[1048][14]);
mul_8x8bit m3146 (image[405],filter[5],mul_out[1048][15]);
mul_8x8bit m3147 (image[431],filter[6],mul_out[1049][13]);
mul_8x8bit m3148 (image[432],filter[7],mul_out[1049][14]);
mul_8x8bit m3149 (image[433],filter[8],mul_out[1049][15]);

adder_8bit ad349 (mul_out[1047][13],mul_out[1047][14],mul_out[1047][15],mul_out[1048][13],mul_out[1048][14],mul_out[1048][15],mul_out[1049][13],mul_out[1049][14],mul_out[1049][15],conv_out[349]);



mul_8x8bit m3150 (image[376],filter[0],mul_out[1050][13]);
mul_8x8bit m3151 (image[377],filter[1],mul_out[1050][14]);
mul_8x8bit m3152 (image[378],filter[2],mul_out[1050][15]);
mul_8x8bit m3153 (image[404],filter[3],mul_out[1051][13]);
mul_8x8bit m3154 (image[405],filter[4],mul_out[1051][14]);
mul_8x8bit m3155 (image[406],filter[5],mul_out[1051][15]);
mul_8x8bit m3156 (image[432],filter[6],mul_out[1052][13]);
mul_8x8bit m3157 (image[433],filter[7],mul_out[1052][14]);
mul_8x8bit m3158 (image[434],filter[8],mul_out[1052][15]);

adder_8bit ad350 (mul_out[1050][13],mul_out[1050][14],mul_out[1050][15],mul_out[1051][13],mul_out[1051][14],mul_out[1051][15],mul_out[1052][13],mul_out[1052][14],mul_out[1052][15],conv_out[350]);



mul_8x8bit m3159 (image[377],filter[0],mul_out[1053][13]);
mul_8x8bit m3160 (image[378],filter[1],mul_out[1053][14]);
mul_8x8bit m3161 (image[379],filter[2],mul_out[1053][15]);
mul_8x8bit m3162 (image[405],filter[3],mul_out[1054][13]);
mul_8x8bit m3163 (image[406],filter[4],mul_out[1054][14]);
mul_8x8bit m3164 (image[407],filter[5],mul_out[1054][15]);
mul_8x8bit m3165 (image[433],filter[6],mul_out[1055][13]);
mul_8x8bit m3166 (image[434],filter[7],mul_out[1055][14]);
mul_8x8bit m3167 (image[435],filter[8],mul_out[1055][15]);

adder_8bit ad351 (mul_out[1053][13],mul_out[1053][14],mul_out[1053][15],mul_out[1054][13],mul_out[1054][14],mul_out[1054][15],mul_out[1055][13],mul_out[1055][14],mul_out[1055][15],conv_out[351]);



mul_8x8bit m3168 (image[378],filter[0],mul_out[1056][13]);
mul_8x8bit m3169 (image[379],filter[1],mul_out[1056][14]);
mul_8x8bit m3170 (image[380],filter[2],mul_out[1056][15]);
mul_8x8bit m3171 (image[406],filter[3],mul_out[1057][13]);
mul_8x8bit m3172 (image[407],filter[4],mul_out[1057][14]);
mul_8x8bit m3173 (image[408],filter[5],mul_out[1057][15]);
mul_8x8bit m3174 (image[434],filter[6],mul_out[1058][13]);
mul_8x8bit m3175 (image[435],filter[7],mul_out[1058][14]);
mul_8x8bit m3176 (image[436],filter[8],mul_out[1058][15]);

adder_8bit ad352 (mul_out[1056][13],mul_out[1056][14],mul_out[1056][15],mul_out[1057][13],mul_out[1057][14],mul_out[1057][15],mul_out[1058][13],mul_out[1058][14],mul_out[1058][15],conv_out[352]);



mul_8x8bit m3177 (image[379],filter[0],mul_out[1059][13]);
mul_8x8bit m3178 (image[380],filter[1],mul_out[1059][14]);
mul_8x8bit m3179 (image[381],filter[2],mul_out[1059][15]);
mul_8x8bit m3180 (image[407],filter[3],mul_out[1060][13]);
mul_8x8bit m3181 (image[408],filter[4],mul_out[1060][14]);
mul_8x8bit m3182 (image[409],filter[5],mul_out[1060][15]);
mul_8x8bit m3183 (image[435],filter[6],mul_out[1061][13]);
mul_8x8bit m3184 (image[436],filter[7],mul_out[1061][14]);
mul_8x8bit m3185 (image[437],filter[8],mul_out[1061][15]);

adder_8bit ad353 (mul_out[1059][13],mul_out[1059][14],mul_out[1059][15],mul_out[1060][13],mul_out[1060][14],mul_out[1060][15],mul_out[1061][13],mul_out[1061][14],mul_out[1061][15],conv_out[353]);



mul_8x8bit m3186 (image[380],filter[0],mul_out[1062][13]);
mul_8x8bit m3187 (image[381],filter[1],mul_out[1062][14]);
mul_8x8bit m3188 (image[382],filter[2],mul_out[1062][15]);
mul_8x8bit m3189 (image[408],filter[3],mul_out[1063][13]);
mul_8x8bit m3190 (image[409],filter[4],mul_out[1063][14]);
mul_8x8bit m3191 (image[410],filter[5],mul_out[1063][15]);
mul_8x8bit m3192 (image[436],filter[6],mul_out[1064][13]);
mul_8x8bit m3193 (image[437],filter[7],mul_out[1064][14]);
mul_8x8bit m3194 (image[438],filter[8],mul_out[1064][15]);

adder_8bit ad354 (mul_out[1062][13],mul_out[1062][14],mul_out[1062][15],mul_out[1063][13],mul_out[1063][14],mul_out[1063][15],mul_out[1064][13],mul_out[1064][14],mul_out[1064][15],conv_out[354]);



mul_8x8bit m3195 (image[381],filter[0],mul_out[1065][13]);
mul_8x8bit m3196 (image[382],filter[1],mul_out[1065][14]);
mul_8x8bit m3197 (image[383],filter[2],mul_out[1065][15]);
mul_8x8bit m3198 (image[409],filter[3],mul_out[1066][13]);
mul_8x8bit m3199 (image[410],filter[4],mul_out[1066][14]);
mul_8x8bit m3200 (image[411],filter[5],mul_out[1066][15]);
mul_8x8bit m3201 (image[437],filter[6],mul_out[1067][13]);
mul_8x8bit m3202 (image[438],filter[7],mul_out[1067][14]);
mul_8x8bit m3203 (image[439],filter[8],mul_out[1067][15]);

adder_8bit ad355 (mul_out[1065][13],mul_out[1065][14],mul_out[1065][15],mul_out[1066][13],mul_out[1066][14],mul_out[1066][15],mul_out[1067][13],mul_out[1067][14],mul_out[1067][15],conv_out[355]);



mul_8x8bit m3204 (image[382],filter[0],mul_out[1068][13]);
mul_8x8bit m3205 (image[383],filter[1],mul_out[1068][14]);
mul_8x8bit m3206 (image[384],filter[2],mul_out[1068][15]);
mul_8x8bit m3207 (image[410],filter[3],mul_out[1069][13]);
mul_8x8bit m3208 (image[411],filter[4],mul_out[1069][14]);
mul_8x8bit m3209 (image[412],filter[5],mul_out[1069][15]);
mul_8x8bit m3210 (image[438],filter[6],mul_out[1070][13]);
mul_8x8bit m3211 (image[439],filter[7],mul_out[1070][14]);
mul_8x8bit m3212 (image[440],filter[8],mul_out[1070][15]);

adder_8bit ad356 (mul_out[1068][13],mul_out[1068][14],mul_out[1068][15],mul_out[1069][13],mul_out[1069][14],mul_out[1069][15],mul_out[1070][13],mul_out[1070][14],mul_out[1070][15],conv_out[356]);



mul_8x8bit m3213 (image[383],filter[0],mul_out[1071][13]);
mul_8x8bit m3214 (image[384],filter[1],mul_out[1071][14]);
mul_8x8bit m3215 (image[385],filter[2],mul_out[1071][15]);
mul_8x8bit m3216 (image[411],filter[3],mul_out[1072][13]);
mul_8x8bit m3217 (image[412],filter[4],mul_out[1072][14]);
mul_8x8bit m3218 (image[413],filter[5],mul_out[1072][15]);
mul_8x8bit m3219 (image[439],filter[6],mul_out[1073][13]);
mul_8x8bit m3220 (image[440],filter[7],mul_out[1073][14]);
mul_8x8bit m3221 (image[441],filter[8],mul_out[1073][15]);

adder_8bit ad357 (mul_out[1071][13],mul_out[1071][14],mul_out[1071][15],mul_out[1072][13],mul_out[1072][14],mul_out[1072][15],mul_out[1073][13],mul_out[1073][14],mul_out[1073][15],conv_out[357]);



mul_8x8bit m3222 (image[384],filter[0],mul_out[1074][13]);
mul_8x8bit m3223 (image[385],filter[1],mul_out[1074][14]);
mul_8x8bit m3224 (image[386],filter[2],mul_out[1074][15]);
mul_8x8bit m3225 (image[412],filter[3],mul_out[1075][13]);
mul_8x8bit m3226 (image[413],filter[4],mul_out[1075][14]);
mul_8x8bit m3227 (image[414],filter[5],mul_out[1075][15]);
mul_8x8bit m3228 (image[440],filter[6],mul_out[1076][13]);
mul_8x8bit m3229 (image[441],filter[7],mul_out[1076][14]);
mul_8x8bit m3230 (image[442],filter[8],mul_out[1076][15]);

adder_8bit ad358 (mul_out[1074][13],mul_out[1074][14],mul_out[1074][15],mul_out[1075][13],mul_out[1075][14],mul_out[1075][15],mul_out[1076][13],mul_out[1076][14],mul_out[1076][15],conv_out[358]);



mul_8x8bit m3231 (image[385],filter[0],mul_out[1077][13]);
mul_8x8bit m3232 (image[386],filter[1],mul_out[1077][14]);
mul_8x8bit m3233 (image[387],filter[2],mul_out[1077][15]);
mul_8x8bit m3234 (image[413],filter[3],mul_out[1078][13]);
mul_8x8bit m3235 (image[414],filter[4],mul_out[1078][14]);
mul_8x8bit m3236 (image[415],filter[5],mul_out[1078][15]);
mul_8x8bit m3237 (image[441],filter[6],mul_out[1079][13]);
mul_8x8bit m3238 (image[442],filter[7],mul_out[1079][14]);
mul_8x8bit m3239 (image[443],filter[8],mul_out[1079][15]);

adder_8bit ad359 (mul_out[1077][13],mul_out[1077][14],mul_out[1077][15],mul_out[1078][13],mul_out[1078][14],mul_out[1078][15],mul_out[1079][13],mul_out[1079][14],mul_out[1079][15],conv_out[359]);



mul_8x8bit m3240 (image[386],filter[0],mul_out[1080][13]);
mul_8x8bit m3241 (image[387],filter[1],mul_out[1080][14]);
mul_8x8bit m3242 (image[388],filter[2],mul_out[1080][15]);
mul_8x8bit m3243 (image[414],filter[3],mul_out[1081][13]);
mul_8x8bit m3244 (image[415],filter[4],mul_out[1081][14]);
mul_8x8bit m3245 (image[416],filter[5],mul_out[1081][15]);
mul_8x8bit m3246 (image[442],filter[6],mul_out[1082][13]);
mul_8x8bit m3247 (image[443],filter[7],mul_out[1082][14]);
mul_8x8bit m3248 (image[444],filter[8],mul_out[1082][15]);

adder_8bit ad360 (mul_out[1080][13],mul_out[1080][14],mul_out[1080][15],mul_out[1081][13],mul_out[1081][14],mul_out[1081][15],mul_out[1082][13],mul_out[1082][14],mul_out[1082][15],conv_out[360]);



mul_8x8bit m3249 (image[387],filter[0],mul_out[1083][13]);
mul_8x8bit m3250 (image[388],filter[1],mul_out[1083][14]);
mul_8x8bit m3251 (image[389],filter[2],mul_out[1083][15]);
mul_8x8bit m3252 (image[415],filter[3],mul_out[1084][13]);
mul_8x8bit m3253 (image[416],filter[4],mul_out[1084][14]);
mul_8x8bit m3254 (image[417],filter[5],mul_out[1084][15]);
mul_8x8bit m3255 (image[443],filter[6],mul_out[1085][13]);
mul_8x8bit m3256 (image[444],filter[7],mul_out[1085][14]);
mul_8x8bit m3257 (image[445],filter[8],mul_out[1085][15]);

adder_8bit ad361 (mul_out[1083][13],mul_out[1083][14],mul_out[1083][15],mul_out[1084][13],mul_out[1084][14],mul_out[1084][15],mul_out[1085][13],mul_out[1085][14],mul_out[1085][15],conv_out[361]);



mul_8x8bit m3258 (image[388],filter[0],mul_out[1086][13]);
mul_8x8bit m3259 (image[389],filter[1],mul_out[1086][14]);
mul_8x8bit m3260 (image[390],filter[2],mul_out[1086][15]);
mul_8x8bit m3261 (image[416],filter[3],mul_out[1087][13]);
mul_8x8bit m3262 (image[417],filter[4],mul_out[1087][14]);
mul_8x8bit m3263 (image[418],filter[5],mul_out[1087][15]);
mul_8x8bit m3264 (image[444],filter[6],mul_out[1088][13]);
mul_8x8bit m3265 (image[445],filter[7],mul_out[1088][14]);
mul_8x8bit m3266 (image[446],filter[8],mul_out[1088][15]);

adder_8bit ad362 (mul_out[1086][13],mul_out[1086][14],mul_out[1086][15],mul_out[1087][13],mul_out[1087][14],mul_out[1087][15],mul_out[1088][13],mul_out[1088][14],mul_out[1088][15],conv_out[362]);



mul_8x8bit m3267 (image[389],filter[0],mul_out[1089][13]);
mul_8x8bit m3268 (image[390],filter[1],mul_out[1089][14]);
mul_8x8bit m3269 (image[391],filter[2],mul_out[1089][15]);
mul_8x8bit m3270 (image[417],filter[3],mul_out[1090][13]);
mul_8x8bit m3271 (image[418],filter[4],mul_out[1090][14]);
mul_8x8bit m3272 (image[419],filter[5],mul_out[1090][15]);
mul_8x8bit m3273 (image[445],filter[6],mul_out[1091][13]);
mul_8x8bit m3274 (image[446],filter[7],mul_out[1091][14]);
mul_8x8bit m3275 (image[447],filter[8],mul_out[1091][15]);

adder_8bit ad363 (mul_out[1089][13],mul_out[1089][14],mul_out[1089][15],mul_out[1090][13],mul_out[1090][14],mul_out[1090][15],mul_out[1091][13],mul_out[1091][14],mul_out[1091][15],conv_out[363]);



mul_8x8bit m3276 (image[392],filter[0],mul_out[1092][14]);
mul_8x8bit m3277 (image[393],filter[1],mul_out[1092][15]);
mul_8x8bit m3278 (image[394],filter[2],mul_out[1092][16]);
mul_8x8bit m3279 (image[420],filter[3],mul_out[1093][14]);
mul_8x8bit m3280 (image[421],filter[4],mul_out[1093][15]);
mul_8x8bit m3281 (image[422],filter[5],mul_out[1093][16]);
mul_8x8bit m3282 (image[448],filter[6],mul_out[1094][14]);
mul_8x8bit m3283 (image[449],filter[7],mul_out[1094][15]);
mul_8x8bit m3284 (image[450],filter[8],mul_out[1094][16]);

adder_8bit ad364 (mul_out[1092][14],mul_out[1092][15],mul_out[1092][16],mul_out[1093][14],mul_out[1093][15],mul_out[1093][16],mul_out[1094][14],mul_out[1094][15],mul_out[1094][16],conv_out[364]);



mul_8x8bit m3285 (image[393],filter[0],mul_out[1095][14]);
mul_8x8bit m3286 (image[394],filter[1],mul_out[1095][15]);
mul_8x8bit m3287 (image[395],filter[2],mul_out[1095][16]);
mul_8x8bit m3288 (image[421],filter[3],mul_out[1096][14]);
mul_8x8bit m3289 (image[422],filter[4],mul_out[1096][15]);
mul_8x8bit m3290 (image[423],filter[5],mul_out[1096][16]);
mul_8x8bit m3291 (image[449],filter[6],mul_out[1097][14]);
mul_8x8bit m3292 (image[450],filter[7],mul_out[1097][15]);
mul_8x8bit m3293 (image[451],filter[8],mul_out[1097][16]);

adder_8bit ad365 (mul_out[1095][14],mul_out[1095][15],mul_out[1095][16],mul_out[1096][14],mul_out[1096][15],mul_out[1096][16],mul_out[1097][14],mul_out[1097][15],mul_out[1097][16],conv_out[365]);



mul_8x8bit m3294 (image[394],filter[0],mul_out[1098][14]);
mul_8x8bit m3295 (image[395],filter[1],mul_out[1098][15]);
mul_8x8bit m3296 (image[396],filter[2],mul_out[1098][16]);
mul_8x8bit m3297 (image[422],filter[3],mul_out[1099][14]);
mul_8x8bit m3298 (image[423],filter[4],mul_out[1099][15]);
mul_8x8bit m3299 (image[424],filter[5],mul_out[1099][16]);
mul_8x8bit m3300 (image[450],filter[6],mul_out[1100][14]);
mul_8x8bit m3301 (image[451],filter[7],mul_out[1100][15]);
mul_8x8bit m3302 (image[452],filter[8],mul_out[1100][16]);

adder_8bit ad366 (mul_out[1098][14],mul_out[1098][15],mul_out[1098][16],mul_out[1099][14],mul_out[1099][15],mul_out[1099][16],mul_out[1100][14],mul_out[1100][15],mul_out[1100][16],conv_out[366]);



mul_8x8bit m3303 (image[395],filter[0],mul_out[1101][14]);
mul_8x8bit m3304 (image[396],filter[1],mul_out[1101][15]);
mul_8x8bit m3305 (image[397],filter[2],mul_out[1101][16]);
mul_8x8bit m3306 (image[423],filter[3],mul_out[1102][14]);
mul_8x8bit m3307 (image[424],filter[4],mul_out[1102][15]);
mul_8x8bit m3308 (image[425],filter[5],mul_out[1102][16]);
mul_8x8bit m3309 (image[451],filter[6],mul_out[1103][14]);
mul_8x8bit m3310 (image[452],filter[7],mul_out[1103][15]);
mul_8x8bit m3311 (image[453],filter[8],mul_out[1103][16]);

adder_8bit ad367 (mul_out[1101][14],mul_out[1101][15],mul_out[1101][16],mul_out[1102][14],mul_out[1102][15],mul_out[1102][16],mul_out[1103][14],mul_out[1103][15],mul_out[1103][16],conv_out[367]);



mul_8x8bit m3312 (image[396],filter[0],mul_out[1104][14]);
mul_8x8bit m3313 (image[397],filter[1],mul_out[1104][15]);
mul_8x8bit m3314 (image[398],filter[2],mul_out[1104][16]);
mul_8x8bit m3315 (image[424],filter[3],mul_out[1105][14]);
mul_8x8bit m3316 (image[425],filter[4],mul_out[1105][15]);
mul_8x8bit m3317 (image[426],filter[5],mul_out[1105][16]);
mul_8x8bit m3318 (image[452],filter[6],mul_out[1106][14]);
mul_8x8bit m3319 (image[453],filter[7],mul_out[1106][15]);
mul_8x8bit m3320 (image[454],filter[8],mul_out[1106][16]);

adder_8bit ad368 (mul_out[1104][14],mul_out[1104][15],mul_out[1104][16],mul_out[1105][14],mul_out[1105][15],mul_out[1105][16],mul_out[1106][14],mul_out[1106][15],mul_out[1106][16],conv_out[368]);



mul_8x8bit m3321 (image[397],filter[0],mul_out[1107][14]);
mul_8x8bit m3322 (image[398],filter[1],mul_out[1107][15]);
mul_8x8bit m3323 (image[399],filter[2],mul_out[1107][16]);
mul_8x8bit m3324 (image[425],filter[3],mul_out[1108][14]);
mul_8x8bit m3325 (image[426],filter[4],mul_out[1108][15]);
mul_8x8bit m3326 (image[427],filter[5],mul_out[1108][16]);
mul_8x8bit m3327 (image[453],filter[6],mul_out[1109][14]);
mul_8x8bit m3328 (image[454],filter[7],mul_out[1109][15]);
mul_8x8bit m3329 (image[455],filter[8],mul_out[1109][16]);

adder_8bit ad369 (mul_out[1107][14],mul_out[1107][15],mul_out[1107][16],mul_out[1108][14],mul_out[1108][15],mul_out[1108][16],mul_out[1109][14],mul_out[1109][15],mul_out[1109][16],conv_out[369]);



mul_8x8bit m3330 (image[398],filter[0],mul_out[1110][14]);
mul_8x8bit m3331 (image[399],filter[1],mul_out[1110][15]);
mul_8x8bit m3332 (image[400],filter[2],mul_out[1110][16]);
mul_8x8bit m3333 (image[426],filter[3],mul_out[1111][14]);
mul_8x8bit m3334 (image[427],filter[4],mul_out[1111][15]);
mul_8x8bit m3335 (image[428],filter[5],mul_out[1111][16]);
mul_8x8bit m3336 (image[454],filter[6],mul_out[1112][14]);
mul_8x8bit m3337 (image[455],filter[7],mul_out[1112][15]);
mul_8x8bit m3338 (image[456],filter[8],mul_out[1112][16]);

adder_8bit ad370 (mul_out[1110][14],mul_out[1110][15],mul_out[1110][16],mul_out[1111][14],mul_out[1111][15],mul_out[1111][16],mul_out[1112][14],mul_out[1112][15],mul_out[1112][16],conv_out[370]);



mul_8x8bit m3339 (image[399],filter[0],mul_out[1113][14]);
mul_8x8bit m3340 (image[400],filter[1],mul_out[1113][15]);
mul_8x8bit m3341 (image[401],filter[2],mul_out[1113][16]);
mul_8x8bit m3342 (image[427],filter[3],mul_out[1114][14]);
mul_8x8bit m3343 (image[428],filter[4],mul_out[1114][15]);
mul_8x8bit m3344 (image[429],filter[5],mul_out[1114][16]);
mul_8x8bit m3345 (image[455],filter[6],mul_out[1115][14]);
mul_8x8bit m3346 (image[456],filter[7],mul_out[1115][15]);
mul_8x8bit m3347 (image[457],filter[8],mul_out[1115][16]);

adder_8bit ad371 (mul_out[1113][14],mul_out[1113][15],mul_out[1113][16],mul_out[1114][14],mul_out[1114][15],mul_out[1114][16],mul_out[1115][14],mul_out[1115][15],mul_out[1115][16],conv_out[371]);



mul_8x8bit m3348 (image[400],filter[0],mul_out[1116][14]);
mul_8x8bit m3349 (image[401],filter[1],mul_out[1116][15]);
mul_8x8bit m3350 (image[402],filter[2],mul_out[1116][16]);
mul_8x8bit m3351 (image[428],filter[3],mul_out[1117][14]);
mul_8x8bit m3352 (image[429],filter[4],mul_out[1117][15]);
mul_8x8bit m3353 (image[430],filter[5],mul_out[1117][16]);
mul_8x8bit m3354 (image[456],filter[6],mul_out[1118][14]);
mul_8x8bit m3355 (image[457],filter[7],mul_out[1118][15]);
mul_8x8bit m3356 (image[458],filter[8],mul_out[1118][16]);

adder_8bit ad372 (mul_out[1116][14],mul_out[1116][15],mul_out[1116][16],mul_out[1117][14],mul_out[1117][15],mul_out[1117][16],mul_out[1118][14],mul_out[1118][15],mul_out[1118][16],conv_out[372]);



mul_8x8bit m3357 (image[401],filter[0],mul_out[1119][14]);
mul_8x8bit m3358 (image[402],filter[1],mul_out[1119][15]);
mul_8x8bit m3359 (image[403],filter[2],mul_out[1119][16]);
mul_8x8bit m3360 (image[429],filter[3],mul_out[1120][14]);
mul_8x8bit m3361 (image[430],filter[4],mul_out[1120][15]);
mul_8x8bit m3362 (image[431],filter[5],mul_out[1120][16]);
mul_8x8bit m3363 (image[457],filter[6],mul_out[1121][14]);
mul_8x8bit m3364 (image[458],filter[7],mul_out[1121][15]);
mul_8x8bit m3365 (image[459],filter[8],mul_out[1121][16]);

adder_8bit ad373 (mul_out[1119][14],mul_out[1119][15],mul_out[1119][16],mul_out[1120][14],mul_out[1120][15],mul_out[1120][16],mul_out[1121][14],mul_out[1121][15],mul_out[1121][16],conv_out[373]);



mul_8x8bit m3366 (image[402],filter[0],mul_out[1122][14]);
mul_8x8bit m3367 (image[403],filter[1],mul_out[1122][15]);
mul_8x8bit m3368 (image[404],filter[2],mul_out[1122][16]);
mul_8x8bit m3369 (image[430],filter[3],mul_out[1123][14]);
mul_8x8bit m3370 (image[431],filter[4],mul_out[1123][15]);
mul_8x8bit m3371 (image[432],filter[5],mul_out[1123][16]);
mul_8x8bit m3372 (image[458],filter[6],mul_out[1124][14]);
mul_8x8bit m3373 (image[459],filter[7],mul_out[1124][15]);
mul_8x8bit m3374 (image[460],filter[8],mul_out[1124][16]);

adder_8bit ad374 (mul_out[1122][14],mul_out[1122][15],mul_out[1122][16],mul_out[1123][14],mul_out[1123][15],mul_out[1123][16],mul_out[1124][14],mul_out[1124][15],mul_out[1124][16],conv_out[374]);



mul_8x8bit m3375 (image[403],filter[0],mul_out[1125][14]);
mul_8x8bit m3376 (image[404],filter[1],mul_out[1125][15]);
mul_8x8bit m3377 (image[405],filter[2],mul_out[1125][16]);
mul_8x8bit m3378 (image[431],filter[3],mul_out[1126][14]);
mul_8x8bit m3379 (image[432],filter[4],mul_out[1126][15]);
mul_8x8bit m3380 (image[433],filter[5],mul_out[1126][16]);
mul_8x8bit m3381 (image[459],filter[6],mul_out[1127][14]);
mul_8x8bit m3382 (image[460],filter[7],mul_out[1127][15]);
mul_8x8bit m3383 (image[461],filter[8],mul_out[1127][16]);

adder_8bit ad375 (mul_out[1125][14],mul_out[1125][15],mul_out[1125][16],mul_out[1126][14],mul_out[1126][15],mul_out[1126][16],mul_out[1127][14],mul_out[1127][15],mul_out[1127][16],conv_out[375]);



mul_8x8bit m3384 (image[404],filter[0],mul_out[1128][14]);
mul_8x8bit m3385 (image[405],filter[1],mul_out[1128][15]);
mul_8x8bit m3386 (image[406],filter[2],mul_out[1128][16]);
mul_8x8bit m3387 (image[432],filter[3],mul_out[1129][14]);
mul_8x8bit m3388 (image[433],filter[4],mul_out[1129][15]);
mul_8x8bit m3389 (image[434],filter[5],mul_out[1129][16]);
mul_8x8bit m3390 (image[460],filter[6],mul_out[1130][14]);
mul_8x8bit m3391 (image[461],filter[7],mul_out[1130][15]);
mul_8x8bit m3392 (image[462],filter[8],mul_out[1130][16]);

adder_8bit ad376 (mul_out[1128][14],mul_out[1128][15],mul_out[1128][16],mul_out[1129][14],mul_out[1129][15],mul_out[1129][16],mul_out[1130][14],mul_out[1130][15],mul_out[1130][16],conv_out[376]);



mul_8x8bit m3393 (image[405],filter[0],mul_out[1131][14]);
mul_8x8bit m3394 (image[406],filter[1],mul_out[1131][15]);
mul_8x8bit m3395 (image[407],filter[2],mul_out[1131][16]);
mul_8x8bit m3396 (image[433],filter[3],mul_out[1132][14]);
mul_8x8bit m3397 (image[434],filter[4],mul_out[1132][15]);
mul_8x8bit m3398 (image[435],filter[5],mul_out[1132][16]);
mul_8x8bit m3399 (image[461],filter[6],mul_out[1133][14]);
mul_8x8bit m3400 (image[462],filter[7],mul_out[1133][15]);
mul_8x8bit m3401 (image[463],filter[8],mul_out[1133][16]);

adder_8bit ad377 (mul_out[1131][14],mul_out[1131][15],mul_out[1131][16],mul_out[1132][14],mul_out[1132][15],mul_out[1132][16],mul_out[1133][14],mul_out[1133][15],mul_out[1133][16],conv_out[377]);



mul_8x8bit m3402 (image[406],filter[0],mul_out[1134][14]);
mul_8x8bit m3403 (image[407],filter[1],mul_out[1134][15]);
mul_8x8bit m3404 (image[408],filter[2],mul_out[1134][16]);
mul_8x8bit m3405 (image[434],filter[3],mul_out[1135][14]);
mul_8x8bit m3406 (image[435],filter[4],mul_out[1135][15]);
mul_8x8bit m3407 (image[436],filter[5],mul_out[1135][16]);
mul_8x8bit m3408 (image[462],filter[6],mul_out[1136][14]);
mul_8x8bit m3409 (image[463],filter[7],mul_out[1136][15]);
mul_8x8bit m3410 (image[464],filter[8],mul_out[1136][16]);

adder_8bit ad378 (mul_out[1134][14],mul_out[1134][15],mul_out[1134][16],mul_out[1135][14],mul_out[1135][15],mul_out[1135][16],mul_out[1136][14],mul_out[1136][15],mul_out[1136][16],conv_out[378]);



mul_8x8bit m3411 (image[407],filter[0],mul_out[1137][14]);
mul_8x8bit m3412 (image[408],filter[1],mul_out[1137][15]);
mul_8x8bit m3413 (image[409],filter[2],mul_out[1137][16]);
mul_8x8bit m3414 (image[435],filter[3],mul_out[1138][14]);
mul_8x8bit m3415 (image[436],filter[4],mul_out[1138][15]);
mul_8x8bit m3416 (image[437],filter[5],mul_out[1138][16]);
mul_8x8bit m3417 (image[463],filter[6],mul_out[1139][14]);
mul_8x8bit m3418 (image[464],filter[7],mul_out[1139][15]);
mul_8x8bit m3419 (image[465],filter[8],mul_out[1139][16]);

adder_8bit ad379 (mul_out[1137][14],mul_out[1137][15],mul_out[1137][16],mul_out[1138][14],mul_out[1138][15],mul_out[1138][16],mul_out[1139][14],mul_out[1139][15],mul_out[1139][16],conv_out[379]);



mul_8x8bit m3420 (image[408],filter[0],mul_out[1140][14]);
mul_8x8bit m3421 (image[409],filter[1],mul_out[1140][15]);
mul_8x8bit m3422 (image[410],filter[2],mul_out[1140][16]);
mul_8x8bit m3423 (image[436],filter[3],mul_out[1141][14]);
mul_8x8bit m3424 (image[437],filter[4],mul_out[1141][15]);
mul_8x8bit m3425 (image[438],filter[5],mul_out[1141][16]);
mul_8x8bit m3426 (image[464],filter[6],mul_out[1142][14]);
mul_8x8bit m3427 (image[465],filter[7],mul_out[1142][15]);
mul_8x8bit m3428 (image[466],filter[8],mul_out[1142][16]);

adder_8bit ad380 (mul_out[1140][14],mul_out[1140][15],mul_out[1140][16],mul_out[1141][14],mul_out[1141][15],mul_out[1141][16],mul_out[1142][14],mul_out[1142][15],mul_out[1142][16],conv_out[380]);



mul_8x8bit m3429 (image[409],filter[0],mul_out[1143][14]);
mul_8x8bit m3430 (image[410],filter[1],mul_out[1143][15]);
mul_8x8bit m3431 (image[411],filter[2],mul_out[1143][16]);
mul_8x8bit m3432 (image[437],filter[3],mul_out[1144][14]);
mul_8x8bit m3433 (image[438],filter[4],mul_out[1144][15]);
mul_8x8bit m3434 (image[439],filter[5],mul_out[1144][16]);
mul_8x8bit m3435 (image[465],filter[6],mul_out[1145][14]);
mul_8x8bit m3436 (image[466],filter[7],mul_out[1145][15]);
mul_8x8bit m3437 (image[467],filter[8],mul_out[1145][16]);

adder_8bit ad381 (mul_out[1143][14],mul_out[1143][15],mul_out[1143][16],mul_out[1144][14],mul_out[1144][15],mul_out[1144][16],mul_out[1145][14],mul_out[1145][15],mul_out[1145][16],conv_out[381]);



mul_8x8bit m3438 (image[410],filter[0],mul_out[1146][14]);
mul_8x8bit m3439 (image[411],filter[1],mul_out[1146][15]);
mul_8x8bit m3440 (image[412],filter[2],mul_out[1146][16]);
mul_8x8bit m3441 (image[438],filter[3],mul_out[1147][14]);
mul_8x8bit m3442 (image[439],filter[4],mul_out[1147][15]);
mul_8x8bit m3443 (image[440],filter[5],mul_out[1147][16]);
mul_8x8bit m3444 (image[466],filter[6],mul_out[1148][14]);
mul_8x8bit m3445 (image[467],filter[7],mul_out[1148][15]);
mul_8x8bit m3446 (image[468],filter[8],mul_out[1148][16]);

adder_8bit ad382 (mul_out[1146][14],mul_out[1146][15],mul_out[1146][16],mul_out[1147][14],mul_out[1147][15],mul_out[1147][16],mul_out[1148][14],mul_out[1148][15],mul_out[1148][16],conv_out[382]);



mul_8x8bit m3447 (image[411],filter[0],mul_out[1149][14]);
mul_8x8bit m3448 (image[412],filter[1],mul_out[1149][15]);
mul_8x8bit m3449 (image[413],filter[2],mul_out[1149][16]);
mul_8x8bit m3450 (image[439],filter[3],mul_out[1150][14]);
mul_8x8bit m3451 (image[440],filter[4],mul_out[1150][15]);
mul_8x8bit m3452 (image[441],filter[5],mul_out[1150][16]);
mul_8x8bit m3453 (image[467],filter[6],mul_out[1151][14]);
mul_8x8bit m3454 (image[468],filter[7],mul_out[1151][15]);
mul_8x8bit m3455 (image[469],filter[8],mul_out[1151][16]);

adder_8bit ad383 (mul_out[1149][14],mul_out[1149][15],mul_out[1149][16],mul_out[1150][14],mul_out[1150][15],mul_out[1150][16],mul_out[1151][14],mul_out[1151][15],mul_out[1151][16],conv_out[383]);



mul_8x8bit m3456 (image[412],filter[0],mul_out[1152][14]);
mul_8x8bit m3457 (image[413],filter[1],mul_out[1152][15]);
mul_8x8bit m3458 (image[414],filter[2],mul_out[1152][16]);
mul_8x8bit m3459 (image[440],filter[3],mul_out[1153][14]);
mul_8x8bit m3460 (image[441],filter[4],mul_out[1153][15]);
mul_8x8bit m3461 (image[442],filter[5],mul_out[1153][16]);
mul_8x8bit m3462 (image[468],filter[6],mul_out[1154][14]);
mul_8x8bit m3463 (image[469],filter[7],mul_out[1154][15]);
mul_8x8bit m3464 (image[470],filter[8],mul_out[1154][16]);

adder_8bit ad384 (mul_out[1152][14],mul_out[1152][15],mul_out[1152][16],mul_out[1153][14],mul_out[1153][15],mul_out[1153][16],mul_out[1154][14],mul_out[1154][15],mul_out[1154][16],conv_out[384]);



mul_8x8bit m3465 (image[413],filter[0],mul_out[1155][14]);
mul_8x8bit m3466 (image[414],filter[1],mul_out[1155][15]);
mul_8x8bit m3467 (image[415],filter[2],mul_out[1155][16]);
mul_8x8bit m3468 (image[441],filter[3],mul_out[1156][14]);
mul_8x8bit m3469 (image[442],filter[4],mul_out[1156][15]);
mul_8x8bit m3470 (image[443],filter[5],mul_out[1156][16]);
mul_8x8bit m3471 (image[469],filter[6],mul_out[1157][14]);
mul_8x8bit m3472 (image[470],filter[7],mul_out[1157][15]);
mul_8x8bit m3473 (image[471],filter[8],mul_out[1157][16]);

adder_8bit ad385 (mul_out[1155][14],mul_out[1155][15],mul_out[1155][16],mul_out[1156][14],mul_out[1156][15],mul_out[1156][16],mul_out[1157][14],mul_out[1157][15],mul_out[1157][16],conv_out[385]);



mul_8x8bit m3474 (image[414],filter[0],mul_out[1158][14]);
mul_8x8bit m3475 (image[415],filter[1],mul_out[1158][15]);
mul_8x8bit m3476 (image[416],filter[2],mul_out[1158][16]);
mul_8x8bit m3477 (image[442],filter[3],mul_out[1159][14]);
mul_8x8bit m3478 (image[443],filter[4],mul_out[1159][15]);
mul_8x8bit m3479 (image[444],filter[5],mul_out[1159][16]);
mul_8x8bit m3480 (image[470],filter[6],mul_out[1160][14]);
mul_8x8bit m3481 (image[471],filter[7],mul_out[1160][15]);
mul_8x8bit m3482 (image[472],filter[8],mul_out[1160][16]);

adder_8bit ad386 (mul_out[1158][14],mul_out[1158][15],mul_out[1158][16],mul_out[1159][14],mul_out[1159][15],mul_out[1159][16],mul_out[1160][14],mul_out[1160][15],mul_out[1160][16],conv_out[386]);



mul_8x8bit m3483 (image[415],filter[0],mul_out[1161][14]);
mul_8x8bit m3484 (image[416],filter[1],mul_out[1161][15]);
mul_8x8bit m3485 (image[417],filter[2],mul_out[1161][16]);
mul_8x8bit m3486 (image[443],filter[3],mul_out[1162][14]);
mul_8x8bit m3487 (image[444],filter[4],mul_out[1162][15]);
mul_8x8bit m3488 (image[445],filter[5],mul_out[1162][16]);
mul_8x8bit m3489 (image[471],filter[6],mul_out[1163][14]);
mul_8x8bit m3490 (image[472],filter[7],mul_out[1163][15]);
mul_8x8bit m3491 (image[473],filter[8],mul_out[1163][16]);

adder_8bit ad387 (mul_out[1161][14],mul_out[1161][15],mul_out[1161][16],mul_out[1162][14],mul_out[1162][15],mul_out[1162][16],mul_out[1163][14],mul_out[1163][15],mul_out[1163][16],conv_out[387]);



mul_8x8bit m3492 (image[416],filter[0],mul_out[1164][14]);
mul_8x8bit m3493 (image[417],filter[1],mul_out[1164][15]);
mul_8x8bit m3494 (image[418],filter[2],mul_out[1164][16]);
mul_8x8bit m3495 (image[444],filter[3],mul_out[1165][14]);
mul_8x8bit m3496 (image[445],filter[4],mul_out[1165][15]);
mul_8x8bit m3497 (image[446],filter[5],mul_out[1165][16]);
mul_8x8bit m3498 (image[472],filter[6],mul_out[1166][14]);
mul_8x8bit m3499 (image[473],filter[7],mul_out[1166][15]);
mul_8x8bit m3500 (image[474],filter[8],mul_out[1166][16]);

adder_8bit ad388 (mul_out[1164][14],mul_out[1164][15],mul_out[1164][16],mul_out[1165][14],mul_out[1165][15],mul_out[1165][16],mul_out[1166][14],mul_out[1166][15],mul_out[1166][16],conv_out[388]);



mul_8x8bit m3501 (image[417],filter[0],mul_out[1167][14]);
mul_8x8bit m3502 (image[418],filter[1],mul_out[1167][15]);
mul_8x8bit m3503 (image[419],filter[2],mul_out[1167][16]);
mul_8x8bit m3504 (image[445],filter[3],mul_out[1168][14]);
mul_8x8bit m3505 (image[446],filter[4],mul_out[1168][15]);
mul_8x8bit m3506 (image[447],filter[5],mul_out[1168][16]);
mul_8x8bit m3507 (image[473],filter[6],mul_out[1169][14]);
mul_8x8bit m3508 (image[474],filter[7],mul_out[1169][15]);
mul_8x8bit m3509 (image[475],filter[8],mul_out[1169][16]);

adder_8bit ad389 (mul_out[1167][14],mul_out[1167][15],mul_out[1167][16],mul_out[1168][14],mul_out[1168][15],mul_out[1168][16],mul_out[1169][14],mul_out[1169][15],mul_out[1169][16],conv_out[389]);



mul_8x8bit m3510 (image[420],filter[0],mul_out[1170][15]);
mul_8x8bit m3511 (image[421],filter[1],mul_out[1170][16]);
mul_8x8bit m3512 (image[422],filter[2],mul_out[1170][17]);
mul_8x8bit m3513 (image[448],filter[3],mul_out[1171][15]);
mul_8x8bit m3514 (image[449],filter[4],mul_out[1171][16]);
mul_8x8bit m3515 (image[450],filter[5],mul_out[1171][17]);
mul_8x8bit m3516 (image[476],filter[6],mul_out[1172][15]);
mul_8x8bit m3517 (image[477],filter[7],mul_out[1172][16]);
mul_8x8bit m3518 (image[478],filter[8],mul_out[1172][17]);

adder_8bit ad390 (mul_out[1170][15],mul_out[1170][16],mul_out[1170][17],mul_out[1171][15],mul_out[1171][16],mul_out[1171][17],mul_out[1172][15],mul_out[1172][16],mul_out[1172][17],conv_out[390]);



mul_8x8bit m3519 (image[421],filter[0],mul_out[1173][15]);
mul_8x8bit m3520 (image[422],filter[1],mul_out[1173][16]);
mul_8x8bit m3521 (image[423],filter[2],mul_out[1173][17]);
mul_8x8bit m3522 (image[449],filter[3],mul_out[1174][15]);
mul_8x8bit m3523 (image[450],filter[4],mul_out[1174][16]);
mul_8x8bit m3524 (image[451],filter[5],mul_out[1174][17]);
mul_8x8bit m3525 (image[477],filter[6],mul_out[1175][15]);
mul_8x8bit m3526 (image[478],filter[7],mul_out[1175][16]);
mul_8x8bit m3527 (image[479],filter[8],mul_out[1175][17]);

adder_8bit ad391 (mul_out[1173][15],mul_out[1173][16],mul_out[1173][17],mul_out[1174][15],mul_out[1174][16],mul_out[1174][17],mul_out[1175][15],mul_out[1175][16],mul_out[1175][17],conv_out[391]);



mul_8x8bit m3528 (image[422],filter[0],mul_out[1176][15]);
mul_8x8bit m3529 (image[423],filter[1],mul_out[1176][16]);
mul_8x8bit m3530 (image[424],filter[2],mul_out[1176][17]);
mul_8x8bit m3531 (image[450],filter[3],mul_out[1177][15]);
mul_8x8bit m3532 (image[451],filter[4],mul_out[1177][16]);
mul_8x8bit m3533 (image[452],filter[5],mul_out[1177][17]);
mul_8x8bit m3534 (image[478],filter[6],mul_out[1178][15]);
mul_8x8bit m3535 (image[479],filter[7],mul_out[1178][16]);
mul_8x8bit m3536 (image[480],filter[8],mul_out[1178][17]);

adder_8bit ad392 (mul_out[1176][15],mul_out[1176][16],mul_out[1176][17],mul_out[1177][15],mul_out[1177][16],mul_out[1177][17],mul_out[1178][15],mul_out[1178][16],mul_out[1178][17],conv_out[392]);



mul_8x8bit m3537 (image[423],filter[0],mul_out[1179][15]);
mul_8x8bit m3538 (image[424],filter[1],mul_out[1179][16]);
mul_8x8bit m3539 (image[425],filter[2],mul_out[1179][17]);
mul_8x8bit m3540 (image[451],filter[3],mul_out[1180][15]);
mul_8x8bit m3541 (image[452],filter[4],mul_out[1180][16]);
mul_8x8bit m3542 (image[453],filter[5],mul_out[1180][17]);
mul_8x8bit m3543 (image[479],filter[6],mul_out[1181][15]);
mul_8x8bit m3544 (image[480],filter[7],mul_out[1181][16]);
mul_8x8bit m3545 (image[481],filter[8],mul_out[1181][17]);

adder_8bit ad393 (mul_out[1179][15],mul_out[1179][16],mul_out[1179][17],mul_out[1180][15],mul_out[1180][16],mul_out[1180][17],mul_out[1181][15],mul_out[1181][16],mul_out[1181][17],conv_out[393]);



mul_8x8bit m3546 (image[424],filter[0],mul_out[1182][15]);
mul_8x8bit m3547 (image[425],filter[1],mul_out[1182][16]);
mul_8x8bit m3548 (image[426],filter[2],mul_out[1182][17]);
mul_8x8bit m3549 (image[452],filter[3],mul_out[1183][15]);
mul_8x8bit m3550 (image[453],filter[4],mul_out[1183][16]);
mul_8x8bit m3551 (image[454],filter[5],mul_out[1183][17]);
mul_8x8bit m3552 (image[480],filter[6],mul_out[1184][15]);
mul_8x8bit m3553 (image[481],filter[7],mul_out[1184][16]);
mul_8x8bit m3554 (image[482],filter[8],mul_out[1184][17]);

adder_8bit ad394 (mul_out[1182][15],mul_out[1182][16],mul_out[1182][17],mul_out[1183][15],mul_out[1183][16],mul_out[1183][17],mul_out[1184][15],mul_out[1184][16],mul_out[1184][17],conv_out[394]);



mul_8x8bit m3555 (image[425],filter[0],mul_out[1185][15]);
mul_8x8bit m3556 (image[426],filter[1],mul_out[1185][16]);
mul_8x8bit m3557 (image[427],filter[2],mul_out[1185][17]);
mul_8x8bit m3558 (image[453],filter[3],mul_out[1186][15]);
mul_8x8bit m3559 (image[454],filter[4],mul_out[1186][16]);
mul_8x8bit m3560 (image[455],filter[5],mul_out[1186][17]);
mul_8x8bit m3561 (image[481],filter[6],mul_out[1187][15]);
mul_8x8bit m3562 (image[482],filter[7],mul_out[1187][16]);
mul_8x8bit m3563 (image[483],filter[8],mul_out[1187][17]);

adder_8bit ad395 (mul_out[1185][15],mul_out[1185][16],mul_out[1185][17],mul_out[1186][15],mul_out[1186][16],mul_out[1186][17],mul_out[1187][15],mul_out[1187][16],mul_out[1187][17],conv_out[395]);



mul_8x8bit m3564 (image[426],filter[0],mul_out[1188][15]);
mul_8x8bit m3565 (image[427],filter[1],mul_out[1188][16]);
mul_8x8bit m3566 (image[428],filter[2],mul_out[1188][17]);
mul_8x8bit m3567 (image[454],filter[3],mul_out[1189][15]);
mul_8x8bit m3568 (image[455],filter[4],mul_out[1189][16]);
mul_8x8bit m3569 (image[456],filter[5],mul_out[1189][17]);
mul_8x8bit m3570 (image[482],filter[6],mul_out[1190][15]);
mul_8x8bit m3571 (image[483],filter[7],mul_out[1190][16]);
mul_8x8bit m3572 (image[484],filter[8],mul_out[1190][17]);

adder_8bit ad396 (mul_out[1188][15],mul_out[1188][16],mul_out[1188][17],mul_out[1189][15],mul_out[1189][16],mul_out[1189][17],mul_out[1190][15],mul_out[1190][16],mul_out[1190][17],conv_out[396]);



mul_8x8bit m3573 (image[427],filter[0],mul_out[1191][15]);
mul_8x8bit m3574 (image[428],filter[1],mul_out[1191][16]);
mul_8x8bit m3575 (image[429],filter[2],mul_out[1191][17]);
mul_8x8bit m3576 (image[455],filter[3],mul_out[1192][15]);
mul_8x8bit m3577 (image[456],filter[4],mul_out[1192][16]);
mul_8x8bit m3578 (image[457],filter[5],mul_out[1192][17]);
mul_8x8bit m3579 (image[483],filter[6],mul_out[1193][15]);
mul_8x8bit m3580 (image[484],filter[7],mul_out[1193][16]);
mul_8x8bit m3581 (image[485],filter[8],mul_out[1193][17]);

adder_8bit ad397 (mul_out[1191][15],mul_out[1191][16],mul_out[1191][17],mul_out[1192][15],mul_out[1192][16],mul_out[1192][17],mul_out[1193][15],mul_out[1193][16],mul_out[1193][17],conv_out[397]);



mul_8x8bit m3582 (image[428],filter[0],mul_out[1194][15]);
mul_8x8bit m3583 (image[429],filter[1],mul_out[1194][16]);
mul_8x8bit m3584 (image[430],filter[2],mul_out[1194][17]);
mul_8x8bit m3585 (image[456],filter[3],mul_out[1195][15]);
mul_8x8bit m3586 (image[457],filter[4],mul_out[1195][16]);
mul_8x8bit m3587 (image[458],filter[5],mul_out[1195][17]);
mul_8x8bit m3588 (image[484],filter[6],mul_out[1196][15]);
mul_8x8bit m3589 (image[485],filter[7],mul_out[1196][16]);
mul_8x8bit m3590 (image[486],filter[8],mul_out[1196][17]);

adder_8bit ad398 (mul_out[1194][15],mul_out[1194][16],mul_out[1194][17],mul_out[1195][15],mul_out[1195][16],mul_out[1195][17],mul_out[1196][15],mul_out[1196][16],mul_out[1196][17],conv_out[398]);



mul_8x8bit m3591 (image[429],filter[0],mul_out[1197][15]);
mul_8x8bit m3592 (image[430],filter[1],mul_out[1197][16]);
mul_8x8bit m3593 (image[431],filter[2],mul_out[1197][17]);
mul_8x8bit m3594 (image[457],filter[3],mul_out[1198][15]);
mul_8x8bit m3595 (image[458],filter[4],mul_out[1198][16]);
mul_8x8bit m3596 (image[459],filter[5],mul_out[1198][17]);
mul_8x8bit m3597 (image[485],filter[6],mul_out[1199][15]);
mul_8x8bit m3598 (image[486],filter[7],mul_out[1199][16]);
mul_8x8bit m3599 (image[487],filter[8],mul_out[1199][17]);

adder_8bit ad399 (mul_out[1197][15],mul_out[1197][16],mul_out[1197][17],mul_out[1198][15],mul_out[1198][16],mul_out[1198][17],mul_out[1199][15],mul_out[1199][16],mul_out[1199][17],conv_out[399]);



mul_8x8bit m3600 (image[430],filter[0],mul_out[1200][15]);
mul_8x8bit m3601 (image[431],filter[1],mul_out[1200][16]);
mul_8x8bit m3602 (image[432],filter[2],mul_out[1200][17]);
mul_8x8bit m3603 (image[458],filter[3],mul_out[1201][15]);
mul_8x8bit m3604 (image[459],filter[4],mul_out[1201][16]);
mul_8x8bit m3605 (image[460],filter[5],mul_out[1201][17]);
mul_8x8bit m3606 (image[486],filter[6],mul_out[1202][15]);
mul_8x8bit m3607 (image[487],filter[7],mul_out[1202][16]);
mul_8x8bit m3608 (image[488],filter[8],mul_out[1202][17]);

adder_8bit ad400 (mul_out[1200][15],mul_out[1200][16],mul_out[1200][17],mul_out[1201][15],mul_out[1201][16],mul_out[1201][17],mul_out[1202][15],mul_out[1202][16],mul_out[1202][17],conv_out[400]);



mul_8x8bit m3609 (image[431],filter[0],mul_out[1203][15]);
mul_8x8bit m3610 (image[432],filter[1],mul_out[1203][16]);
mul_8x8bit m3611 (image[433],filter[2],mul_out[1203][17]);
mul_8x8bit m3612 (image[459],filter[3],mul_out[1204][15]);
mul_8x8bit m3613 (image[460],filter[4],mul_out[1204][16]);
mul_8x8bit m3614 (image[461],filter[5],mul_out[1204][17]);
mul_8x8bit m3615 (image[487],filter[6],mul_out[1205][15]);
mul_8x8bit m3616 (image[488],filter[7],mul_out[1205][16]);
mul_8x8bit m3617 (image[489],filter[8],mul_out[1205][17]);

adder_8bit ad401 (mul_out[1203][15],mul_out[1203][16],mul_out[1203][17],mul_out[1204][15],mul_out[1204][16],mul_out[1204][17],mul_out[1205][15],mul_out[1205][16],mul_out[1205][17],conv_out[401]);



mul_8x8bit m3618 (image[432],filter[0],mul_out[1206][15]);
mul_8x8bit m3619 (image[433],filter[1],mul_out[1206][16]);
mul_8x8bit m3620 (image[434],filter[2],mul_out[1206][17]);
mul_8x8bit m3621 (image[460],filter[3],mul_out[1207][15]);
mul_8x8bit m3622 (image[461],filter[4],mul_out[1207][16]);
mul_8x8bit m3623 (image[462],filter[5],mul_out[1207][17]);
mul_8x8bit m3624 (image[488],filter[6],mul_out[1208][15]);
mul_8x8bit m3625 (image[489],filter[7],mul_out[1208][16]);
mul_8x8bit m3626 (image[490],filter[8],mul_out[1208][17]);

adder_8bit ad402 (mul_out[1206][15],mul_out[1206][16],mul_out[1206][17],mul_out[1207][15],mul_out[1207][16],mul_out[1207][17],mul_out[1208][15],mul_out[1208][16],mul_out[1208][17],conv_out[402]);



mul_8x8bit m3627 (image[433],filter[0],mul_out[1209][15]);
mul_8x8bit m3628 (image[434],filter[1],mul_out[1209][16]);
mul_8x8bit m3629 (image[435],filter[2],mul_out[1209][17]);
mul_8x8bit m3630 (image[461],filter[3],mul_out[1210][15]);
mul_8x8bit m3631 (image[462],filter[4],mul_out[1210][16]);
mul_8x8bit m3632 (image[463],filter[5],mul_out[1210][17]);
mul_8x8bit m3633 (image[489],filter[6],mul_out[1211][15]);
mul_8x8bit m3634 (image[490],filter[7],mul_out[1211][16]);
mul_8x8bit m3635 (image[491],filter[8],mul_out[1211][17]);

adder_8bit ad403 (mul_out[1209][15],mul_out[1209][16],mul_out[1209][17],mul_out[1210][15],mul_out[1210][16],mul_out[1210][17],mul_out[1211][15],mul_out[1211][16],mul_out[1211][17],conv_out[403]);



mul_8x8bit m3636 (image[434],filter[0],mul_out[1212][15]);
mul_8x8bit m3637 (image[435],filter[1],mul_out[1212][16]);
mul_8x8bit m3638 (image[436],filter[2],mul_out[1212][17]);
mul_8x8bit m3639 (image[462],filter[3],mul_out[1213][15]);
mul_8x8bit m3640 (image[463],filter[4],mul_out[1213][16]);
mul_8x8bit m3641 (image[464],filter[5],mul_out[1213][17]);
mul_8x8bit m3642 (image[490],filter[6],mul_out[1214][15]);
mul_8x8bit m3643 (image[491],filter[7],mul_out[1214][16]);
mul_8x8bit m3644 (image[492],filter[8],mul_out[1214][17]);

adder_8bit ad404 (mul_out[1212][15],mul_out[1212][16],mul_out[1212][17],mul_out[1213][15],mul_out[1213][16],mul_out[1213][17],mul_out[1214][15],mul_out[1214][16],mul_out[1214][17],conv_out[404]);



mul_8x8bit m3645 (image[435],filter[0],mul_out[1215][15]);
mul_8x8bit m3646 (image[436],filter[1],mul_out[1215][16]);
mul_8x8bit m3647 (image[437],filter[2],mul_out[1215][17]);
mul_8x8bit m3648 (image[463],filter[3],mul_out[1216][15]);
mul_8x8bit m3649 (image[464],filter[4],mul_out[1216][16]);
mul_8x8bit m3650 (image[465],filter[5],mul_out[1216][17]);
mul_8x8bit m3651 (image[491],filter[6],mul_out[1217][15]);
mul_8x8bit m3652 (image[492],filter[7],mul_out[1217][16]);
mul_8x8bit m3653 (image[493],filter[8],mul_out[1217][17]);

adder_8bit ad405 (mul_out[1215][15],mul_out[1215][16],mul_out[1215][17],mul_out[1216][15],mul_out[1216][16],mul_out[1216][17],mul_out[1217][15],mul_out[1217][16],mul_out[1217][17],conv_out[405]);



mul_8x8bit m3654 (image[436],filter[0],mul_out[1218][15]);
mul_8x8bit m3655 (image[437],filter[1],mul_out[1218][16]);
mul_8x8bit m3656 (image[438],filter[2],mul_out[1218][17]);
mul_8x8bit m3657 (image[464],filter[3],mul_out[1219][15]);
mul_8x8bit m3658 (image[465],filter[4],mul_out[1219][16]);
mul_8x8bit m3659 (image[466],filter[5],mul_out[1219][17]);
mul_8x8bit m3660 (image[492],filter[6],mul_out[1220][15]);
mul_8x8bit m3661 (image[493],filter[7],mul_out[1220][16]);
mul_8x8bit m3662 (image[494],filter[8],mul_out[1220][17]);

adder_8bit ad406 (mul_out[1218][15],mul_out[1218][16],mul_out[1218][17],mul_out[1219][15],mul_out[1219][16],mul_out[1219][17],mul_out[1220][15],mul_out[1220][16],mul_out[1220][17],conv_out[406]);



mul_8x8bit m3663 (image[437],filter[0],mul_out[1221][15]);
mul_8x8bit m3664 (image[438],filter[1],mul_out[1221][16]);
mul_8x8bit m3665 (image[439],filter[2],mul_out[1221][17]);
mul_8x8bit m3666 (image[465],filter[3],mul_out[1222][15]);
mul_8x8bit m3667 (image[466],filter[4],mul_out[1222][16]);
mul_8x8bit m3668 (image[467],filter[5],mul_out[1222][17]);
mul_8x8bit m3669 (image[493],filter[6],mul_out[1223][15]);
mul_8x8bit m3670 (image[494],filter[7],mul_out[1223][16]);
mul_8x8bit m3671 (image[495],filter[8],mul_out[1223][17]);

adder_8bit ad407 (mul_out[1221][15],mul_out[1221][16],mul_out[1221][17],mul_out[1222][15],mul_out[1222][16],mul_out[1222][17],mul_out[1223][15],mul_out[1223][16],mul_out[1223][17],conv_out[407]);



mul_8x8bit m3672 (image[438],filter[0],mul_out[1224][15]);
mul_8x8bit m3673 (image[439],filter[1],mul_out[1224][16]);
mul_8x8bit m3674 (image[440],filter[2],mul_out[1224][17]);
mul_8x8bit m3675 (image[466],filter[3],mul_out[1225][15]);
mul_8x8bit m3676 (image[467],filter[4],mul_out[1225][16]);
mul_8x8bit m3677 (image[468],filter[5],mul_out[1225][17]);
mul_8x8bit m3678 (image[494],filter[6],mul_out[1226][15]);
mul_8x8bit m3679 (image[495],filter[7],mul_out[1226][16]);
mul_8x8bit m3680 (image[496],filter[8],mul_out[1226][17]);

adder_8bit ad408 (mul_out[1224][15],mul_out[1224][16],mul_out[1224][17],mul_out[1225][15],mul_out[1225][16],mul_out[1225][17],mul_out[1226][15],mul_out[1226][16],mul_out[1226][17],conv_out[408]);



mul_8x8bit m3681 (image[439],filter[0],mul_out[1227][15]);
mul_8x8bit m3682 (image[440],filter[1],mul_out[1227][16]);
mul_8x8bit m3683 (image[441],filter[2],mul_out[1227][17]);
mul_8x8bit m3684 (image[467],filter[3],mul_out[1228][15]);
mul_8x8bit m3685 (image[468],filter[4],mul_out[1228][16]);
mul_8x8bit m3686 (image[469],filter[5],mul_out[1228][17]);
mul_8x8bit m3687 (image[495],filter[6],mul_out[1229][15]);
mul_8x8bit m3688 (image[496],filter[7],mul_out[1229][16]);
mul_8x8bit m3689 (image[497],filter[8],mul_out[1229][17]);

adder_8bit ad409 (mul_out[1227][15],mul_out[1227][16],mul_out[1227][17],mul_out[1228][15],mul_out[1228][16],mul_out[1228][17],mul_out[1229][15],mul_out[1229][16],mul_out[1229][17],conv_out[409]);



mul_8x8bit m3690 (image[440],filter[0],mul_out[1230][15]);
mul_8x8bit m3691 (image[441],filter[1],mul_out[1230][16]);
mul_8x8bit m3692 (image[442],filter[2],mul_out[1230][17]);
mul_8x8bit m3693 (image[468],filter[3],mul_out[1231][15]);
mul_8x8bit m3694 (image[469],filter[4],mul_out[1231][16]);
mul_8x8bit m3695 (image[470],filter[5],mul_out[1231][17]);
mul_8x8bit m3696 (image[496],filter[6],mul_out[1232][15]);
mul_8x8bit m3697 (image[497],filter[7],mul_out[1232][16]);
mul_8x8bit m3698 (image[498],filter[8],mul_out[1232][17]);

adder_8bit ad410 (mul_out[1230][15],mul_out[1230][16],mul_out[1230][17],mul_out[1231][15],mul_out[1231][16],mul_out[1231][17],mul_out[1232][15],mul_out[1232][16],mul_out[1232][17],conv_out[410]);



mul_8x8bit m3699 (image[441],filter[0],mul_out[1233][15]);
mul_8x8bit m3700 (image[442],filter[1],mul_out[1233][16]);
mul_8x8bit m3701 (image[443],filter[2],mul_out[1233][17]);
mul_8x8bit m3702 (image[469],filter[3],mul_out[1234][15]);
mul_8x8bit m3703 (image[470],filter[4],mul_out[1234][16]);
mul_8x8bit m3704 (image[471],filter[5],mul_out[1234][17]);
mul_8x8bit m3705 (image[497],filter[6],mul_out[1235][15]);
mul_8x8bit m3706 (image[498],filter[7],mul_out[1235][16]);
mul_8x8bit m3707 (image[499],filter[8],mul_out[1235][17]);

adder_8bit ad411 (mul_out[1233][15],mul_out[1233][16],mul_out[1233][17],mul_out[1234][15],mul_out[1234][16],mul_out[1234][17],mul_out[1235][15],mul_out[1235][16],mul_out[1235][17],conv_out[411]);



mul_8x8bit m3708 (image[442],filter[0],mul_out[1236][15]);
mul_8x8bit m3709 (image[443],filter[1],mul_out[1236][16]);
mul_8x8bit m3710 (image[444],filter[2],mul_out[1236][17]);
mul_8x8bit m3711 (image[470],filter[3],mul_out[1237][15]);
mul_8x8bit m3712 (image[471],filter[4],mul_out[1237][16]);
mul_8x8bit m3713 (image[472],filter[5],mul_out[1237][17]);
mul_8x8bit m3714 (image[498],filter[6],mul_out[1238][15]);
mul_8x8bit m3715 (image[499],filter[7],mul_out[1238][16]);
mul_8x8bit m3716 (image[500],filter[8],mul_out[1238][17]);

adder_8bit ad412 (mul_out[1236][15],mul_out[1236][16],mul_out[1236][17],mul_out[1237][15],mul_out[1237][16],mul_out[1237][17],mul_out[1238][15],mul_out[1238][16],mul_out[1238][17],conv_out[412]);



mul_8x8bit m3717 (image[443],filter[0],mul_out[1239][15]);
mul_8x8bit m3718 (image[444],filter[1],mul_out[1239][16]);
mul_8x8bit m3719 (image[445],filter[2],mul_out[1239][17]);
mul_8x8bit m3720 (image[471],filter[3],mul_out[1240][15]);
mul_8x8bit m3721 (image[472],filter[4],mul_out[1240][16]);
mul_8x8bit m3722 (image[473],filter[5],mul_out[1240][17]);
mul_8x8bit m3723 (image[499],filter[6],mul_out[1241][15]);
mul_8x8bit m3724 (image[500],filter[7],mul_out[1241][16]);
mul_8x8bit m3725 (image[501],filter[8],mul_out[1241][17]);

adder_8bit ad413 (mul_out[1239][15],mul_out[1239][16],mul_out[1239][17],mul_out[1240][15],mul_out[1240][16],mul_out[1240][17],mul_out[1241][15],mul_out[1241][16],mul_out[1241][17],conv_out[413]);



mul_8x8bit m3726 (image[444],filter[0],mul_out[1242][15]);
mul_8x8bit m3727 (image[445],filter[1],mul_out[1242][16]);
mul_8x8bit m3728 (image[446],filter[2],mul_out[1242][17]);
mul_8x8bit m3729 (image[472],filter[3],mul_out[1243][15]);
mul_8x8bit m3730 (image[473],filter[4],mul_out[1243][16]);
mul_8x8bit m3731 (image[474],filter[5],mul_out[1243][17]);
mul_8x8bit m3732 (image[500],filter[6],mul_out[1244][15]);
mul_8x8bit m3733 (image[501],filter[7],mul_out[1244][16]);
mul_8x8bit m3734 (image[502],filter[8],mul_out[1244][17]);

adder_8bit ad414 (mul_out[1242][15],mul_out[1242][16],mul_out[1242][17],mul_out[1243][15],mul_out[1243][16],mul_out[1243][17],mul_out[1244][15],mul_out[1244][16],mul_out[1244][17],conv_out[414]);



mul_8x8bit m3735 (image[445],filter[0],mul_out[1245][15]);
mul_8x8bit m3736 (image[446],filter[1],mul_out[1245][16]);
mul_8x8bit m3737 (image[447],filter[2],mul_out[1245][17]);
mul_8x8bit m3738 (image[473],filter[3],mul_out[1246][15]);
mul_8x8bit m3739 (image[474],filter[4],mul_out[1246][16]);
mul_8x8bit m3740 (image[475],filter[5],mul_out[1246][17]);
mul_8x8bit m3741 (image[501],filter[6],mul_out[1247][15]);
mul_8x8bit m3742 (image[502],filter[7],mul_out[1247][16]);
mul_8x8bit m3743 (image[503],filter[8],mul_out[1247][17]);

adder_8bit ad415 (mul_out[1245][15],mul_out[1245][16],mul_out[1245][17],mul_out[1246][15],mul_out[1246][16],mul_out[1246][17],mul_out[1247][15],mul_out[1247][16],mul_out[1247][17],conv_out[415]);



mul_8x8bit m3744 (image[448],filter[0],mul_out[1248][16]);
mul_8x8bit m3745 (image[449],filter[1],mul_out[1248][17]);
mul_8x8bit m3746 (image[450],filter[2],mul_out[1248][18]);
mul_8x8bit m3747 (image[476],filter[3],mul_out[1249][16]);
mul_8x8bit m3748 (image[477],filter[4],mul_out[1249][17]);
mul_8x8bit m3749 (image[478],filter[5],mul_out[1249][18]);
mul_8x8bit m3750 (image[504],filter[6],mul_out[1250][16]);
mul_8x8bit m3751 (image[505],filter[7],mul_out[1250][17]);
mul_8x8bit m3752 (image[506],filter[8],mul_out[1250][18]);

adder_8bit ad416 (mul_out[1248][16],mul_out[1248][17],mul_out[1248][18],mul_out[1249][16],mul_out[1249][17],mul_out[1249][18],mul_out[1250][16],mul_out[1250][17],mul_out[1250][18],conv_out[416]);



mul_8x8bit m3753 (image[449],filter[0],mul_out[1251][16]);
mul_8x8bit m3754 (image[450],filter[1],mul_out[1251][17]);
mul_8x8bit m3755 (image[451],filter[2],mul_out[1251][18]);
mul_8x8bit m3756 (image[477],filter[3],mul_out[1252][16]);
mul_8x8bit m3757 (image[478],filter[4],mul_out[1252][17]);
mul_8x8bit m3758 (image[479],filter[5],mul_out[1252][18]);
mul_8x8bit m3759 (image[505],filter[6],mul_out[1253][16]);
mul_8x8bit m3760 (image[506],filter[7],mul_out[1253][17]);
mul_8x8bit m3761 (image[507],filter[8],mul_out[1253][18]);

adder_8bit ad417 (mul_out[1251][16],mul_out[1251][17],mul_out[1251][18],mul_out[1252][16],mul_out[1252][17],mul_out[1252][18],mul_out[1253][16],mul_out[1253][17],mul_out[1253][18],conv_out[417]);



mul_8x8bit m3762 (image[450],filter[0],mul_out[1254][16]);
mul_8x8bit m3763 (image[451],filter[1],mul_out[1254][17]);
mul_8x8bit m3764 (image[452],filter[2],mul_out[1254][18]);
mul_8x8bit m3765 (image[478],filter[3],mul_out[1255][16]);
mul_8x8bit m3766 (image[479],filter[4],mul_out[1255][17]);
mul_8x8bit m3767 (image[480],filter[5],mul_out[1255][18]);
mul_8x8bit m3768 (image[506],filter[6],mul_out[1256][16]);
mul_8x8bit m3769 (image[507],filter[7],mul_out[1256][17]);
mul_8x8bit m3770 (image[508],filter[8],mul_out[1256][18]);

adder_8bit ad418 (mul_out[1254][16],mul_out[1254][17],mul_out[1254][18],mul_out[1255][16],mul_out[1255][17],mul_out[1255][18],mul_out[1256][16],mul_out[1256][17],mul_out[1256][18],conv_out[418]);



mul_8x8bit m3771 (image[451],filter[0],mul_out[1257][16]);
mul_8x8bit m3772 (image[452],filter[1],mul_out[1257][17]);
mul_8x8bit m3773 (image[453],filter[2],mul_out[1257][18]);
mul_8x8bit m3774 (image[479],filter[3],mul_out[1258][16]);
mul_8x8bit m3775 (image[480],filter[4],mul_out[1258][17]);
mul_8x8bit m3776 (image[481],filter[5],mul_out[1258][18]);
mul_8x8bit m3777 (image[507],filter[6],mul_out[1259][16]);
mul_8x8bit m3778 (image[508],filter[7],mul_out[1259][17]);
mul_8x8bit m3779 (image[509],filter[8],mul_out[1259][18]);

adder_8bit ad419 (mul_out[1257][16],mul_out[1257][17],mul_out[1257][18],mul_out[1258][16],mul_out[1258][17],mul_out[1258][18],mul_out[1259][16],mul_out[1259][17],mul_out[1259][18],conv_out[419]);



mul_8x8bit m3780 (image[452],filter[0],mul_out[1260][16]);
mul_8x8bit m3781 (image[453],filter[1],mul_out[1260][17]);
mul_8x8bit m3782 (image[454],filter[2],mul_out[1260][18]);
mul_8x8bit m3783 (image[480],filter[3],mul_out[1261][16]);
mul_8x8bit m3784 (image[481],filter[4],mul_out[1261][17]);
mul_8x8bit m3785 (image[482],filter[5],mul_out[1261][18]);
mul_8x8bit m3786 (image[508],filter[6],mul_out[1262][16]);
mul_8x8bit m3787 (image[509],filter[7],mul_out[1262][17]);
mul_8x8bit m3788 (image[510],filter[8],mul_out[1262][18]);

adder_8bit ad420 (mul_out[1260][16],mul_out[1260][17],mul_out[1260][18],mul_out[1261][16],mul_out[1261][17],mul_out[1261][18],mul_out[1262][16],mul_out[1262][17],mul_out[1262][18],conv_out[420]);



mul_8x8bit m3789 (image[453],filter[0],mul_out[1263][16]);
mul_8x8bit m3790 (image[454],filter[1],mul_out[1263][17]);
mul_8x8bit m3791 (image[455],filter[2],mul_out[1263][18]);
mul_8x8bit m3792 (image[481],filter[3],mul_out[1264][16]);
mul_8x8bit m3793 (image[482],filter[4],mul_out[1264][17]);
mul_8x8bit m3794 (image[483],filter[5],mul_out[1264][18]);
mul_8x8bit m3795 (image[509],filter[6],mul_out[1265][16]);
mul_8x8bit m3796 (image[510],filter[7],mul_out[1265][17]);
mul_8x8bit m3797 (image[511],filter[8],mul_out[1265][18]);

adder_8bit ad421 (mul_out[1263][16],mul_out[1263][17],mul_out[1263][18],mul_out[1264][16],mul_out[1264][17],mul_out[1264][18],mul_out[1265][16],mul_out[1265][17],mul_out[1265][18],conv_out[421]);



mul_8x8bit m3798 (image[454],filter[0],mul_out[1266][16]);
mul_8x8bit m3799 (image[455],filter[1],mul_out[1266][17]);
mul_8x8bit m3800 (image[456],filter[2],mul_out[1266][18]);
mul_8x8bit m3801 (image[482],filter[3],mul_out[1267][16]);
mul_8x8bit m3802 (image[483],filter[4],mul_out[1267][17]);
mul_8x8bit m3803 (image[484],filter[5],mul_out[1267][18]);
mul_8x8bit m3804 (image[510],filter[6],mul_out[1268][16]);
mul_8x8bit m3805 (image[511],filter[7],mul_out[1268][17]);
mul_8x8bit m3806 (image[512],filter[8],mul_out[1268][18]);

adder_8bit ad422 (mul_out[1266][16],mul_out[1266][17],mul_out[1266][18],mul_out[1267][16],mul_out[1267][17],mul_out[1267][18],mul_out[1268][16],mul_out[1268][17],mul_out[1268][18],conv_out[422]);



mul_8x8bit m3807 (image[455],filter[0],mul_out[1269][16]);
mul_8x8bit m3808 (image[456],filter[1],mul_out[1269][17]);
mul_8x8bit m3809 (image[457],filter[2],mul_out[1269][18]);
mul_8x8bit m3810 (image[483],filter[3],mul_out[1270][16]);
mul_8x8bit m3811 (image[484],filter[4],mul_out[1270][17]);
mul_8x8bit m3812 (image[485],filter[5],mul_out[1270][18]);
mul_8x8bit m3813 (image[511],filter[6],mul_out[1271][16]);
mul_8x8bit m3814 (image[512],filter[7],mul_out[1271][17]);
mul_8x8bit m3815 (image[513],filter[8],mul_out[1271][18]);

adder_8bit ad423 (mul_out[1269][16],mul_out[1269][17],mul_out[1269][18],mul_out[1270][16],mul_out[1270][17],mul_out[1270][18],mul_out[1271][16],mul_out[1271][17],mul_out[1271][18],conv_out[423]);



mul_8x8bit m3816 (image[456],filter[0],mul_out[1272][16]);
mul_8x8bit m3817 (image[457],filter[1],mul_out[1272][17]);
mul_8x8bit m3818 (image[458],filter[2],mul_out[1272][18]);
mul_8x8bit m3819 (image[484],filter[3],mul_out[1273][16]);
mul_8x8bit m3820 (image[485],filter[4],mul_out[1273][17]);
mul_8x8bit m3821 (image[486],filter[5],mul_out[1273][18]);
mul_8x8bit m3822 (image[512],filter[6],mul_out[1274][16]);
mul_8x8bit m3823 (image[513],filter[7],mul_out[1274][17]);
mul_8x8bit m3824 (image[514],filter[8],mul_out[1274][18]);

adder_8bit ad424 (mul_out[1272][16],mul_out[1272][17],mul_out[1272][18],mul_out[1273][16],mul_out[1273][17],mul_out[1273][18],mul_out[1274][16],mul_out[1274][17],mul_out[1274][18],conv_out[424]);



mul_8x8bit m3825 (image[457],filter[0],mul_out[1275][16]);
mul_8x8bit m3826 (image[458],filter[1],mul_out[1275][17]);
mul_8x8bit m3827 (image[459],filter[2],mul_out[1275][18]);
mul_8x8bit m3828 (image[485],filter[3],mul_out[1276][16]);
mul_8x8bit m3829 (image[486],filter[4],mul_out[1276][17]);
mul_8x8bit m3830 (image[487],filter[5],mul_out[1276][18]);
mul_8x8bit m3831 (image[513],filter[6],mul_out[1277][16]);
mul_8x8bit m3832 (image[514],filter[7],mul_out[1277][17]);
mul_8x8bit m3833 (image[515],filter[8],mul_out[1277][18]);

adder_8bit ad425 (mul_out[1275][16],mul_out[1275][17],mul_out[1275][18],mul_out[1276][16],mul_out[1276][17],mul_out[1276][18],mul_out[1277][16],mul_out[1277][17],mul_out[1277][18],conv_out[425]);



mul_8x8bit m3834 (image[458],filter[0],mul_out[1278][16]);
mul_8x8bit m3835 (image[459],filter[1],mul_out[1278][17]);
mul_8x8bit m3836 (image[460],filter[2],mul_out[1278][18]);
mul_8x8bit m3837 (image[486],filter[3],mul_out[1279][16]);
mul_8x8bit m3838 (image[487],filter[4],mul_out[1279][17]);
mul_8x8bit m3839 (image[488],filter[5],mul_out[1279][18]);
mul_8x8bit m3840 (image[514],filter[6],mul_out[1280][16]);
mul_8x8bit m3841 (image[515],filter[7],mul_out[1280][17]);
mul_8x8bit m3842 (image[516],filter[8],mul_out[1280][18]);

adder_8bit ad426 (mul_out[1278][16],mul_out[1278][17],mul_out[1278][18],mul_out[1279][16],mul_out[1279][17],mul_out[1279][18],mul_out[1280][16],mul_out[1280][17],mul_out[1280][18],conv_out[426]);



mul_8x8bit m3843 (image[459],filter[0],mul_out[1281][16]);
mul_8x8bit m3844 (image[460],filter[1],mul_out[1281][17]);
mul_8x8bit m3845 (image[461],filter[2],mul_out[1281][18]);
mul_8x8bit m3846 (image[487],filter[3],mul_out[1282][16]);
mul_8x8bit m3847 (image[488],filter[4],mul_out[1282][17]);
mul_8x8bit m3848 (image[489],filter[5],mul_out[1282][18]);
mul_8x8bit m3849 (image[515],filter[6],mul_out[1283][16]);
mul_8x8bit m3850 (image[516],filter[7],mul_out[1283][17]);
mul_8x8bit m3851 (image[517],filter[8],mul_out[1283][18]);

adder_8bit ad427 (mul_out[1281][16],mul_out[1281][17],mul_out[1281][18],mul_out[1282][16],mul_out[1282][17],mul_out[1282][18],mul_out[1283][16],mul_out[1283][17],mul_out[1283][18],conv_out[427]);



mul_8x8bit m3852 (image[460],filter[0],mul_out[1284][16]);
mul_8x8bit m3853 (image[461],filter[1],mul_out[1284][17]);
mul_8x8bit m3854 (image[462],filter[2],mul_out[1284][18]);
mul_8x8bit m3855 (image[488],filter[3],mul_out[1285][16]);
mul_8x8bit m3856 (image[489],filter[4],mul_out[1285][17]);
mul_8x8bit m3857 (image[490],filter[5],mul_out[1285][18]);
mul_8x8bit m3858 (image[516],filter[6],mul_out[1286][16]);
mul_8x8bit m3859 (image[517],filter[7],mul_out[1286][17]);
mul_8x8bit m3860 (image[518],filter[8],mul_out[1286][18]);

adder_8bit ad428 (mul_out[1284][16],mul_out[1284][17],mul_out[1284][18],mul_out[1285][16],mul_out[1285][17],mul_out[1285][18],mul_out[1286][16],mul_out[1286][17],mul_out[1286][18],conv_out[428]);



mul_8x8bit m3861 (image[461],filter[0],mul_out[1287][16]);
mul_8x8bit m3862 (image[462],filter[1],mul_out[1287][17]);
mul_8x8bit m3863 (image[463],filter[2],mul_out[1287][18]);
mul_8x8bit m3864 (image[489],filter[3],mul_out[1288][16]);
mul_8x8bit m3865 (image[490],filter[4],mul_out[1288][17]);
mul_8x8bit m3866 (image[491],filter[5],mul_out[1288][18]);
mul_8x8bit m3867 (image[517],filter[6],mul_out[1289][16]);
mul_8x8bit m3868 (image[518],filter[7],mul_out[1289][17]);
mul_8x8bit m3869 (image[519],filter[8],mul_out[1289][18]);

adder_8bit ad429 (mul_out[1287][16],mul_out[1287][17],mul_out[1287][18],mul_out[1288][16],mul_out[1288][17],mul_out[1288][18],mul_out[1289][16],mul_out[1289][17],mul_out[1289][18],conv_out[429]);



mul_8x8bit m3870 (image[462],filter[0],mul_out[1290][16]);
mul_8x8bit m3871 (image[463],filter[1],mul_out[1290][17]);
mul_8x8bit m3872 (image[464],filter[2],mul_out[1290][18]);
mul_8x8bit m3873 (image[490],filter[3],mul_out[1291][16]);
mul_8x8bit m3874 (image[491],filter[4],mul_out[1291][17]);
mul_8x8bit m3875 (image[492],filter[5],mul_out[1291][18]);
mul_8x8bit m3876 (image[518],filter[6],mul_out[1292][16]);
mul_8x8bit m3877 (image[519],filter[7],mul_out[1292][17]);
mul_8x8bit m3878 (image[520],filter[8],mul_out[1292][18]);

adder_8bit ad430 (mul_out[1290][16],mul_out[1290][17],mul_out[1290][18],mul_out[1291][16],mul_out[1291][17],mul_out[1291][18],mul_out[1292][16],mul_out[1292][17],mul_out[1292][18],conv_out[430]);



mul_8x8bit m3879 (image[463],filter[0],mul_out[1293][16]);
mul_8x8bit m3880 (image[464],filter[1],mul_out[1293][17]);
mul_8x8bit m3881 (image[465],filter[2],mul_out[1293][18]);
mul_8x8bit m3882 (image[491],filter[3],mul_out[1294][16]);
mul_8x8bit m3883 (image[492],filter[4],mul_out[1294][17]);
mul_8x8bit m3884 (image[493],filter[5],mul_out[1294][18]);
mul_8x8bit m3885 (image[519],filter[6],mul_out[1295][16]);
mul_8x8bit m3886 (image[520],filter[7],mul_out[1295][17]);
mul_8x8bit m3887 (image[521],filter[8],mul_out[1295][18]);

adder_8bit ad431 (mul_out[1293][16],mul_out[1293][17],mul_out[1293][18],mul_out[1294][16],mul_out[1294][17],mul_out[1294][18],mul_out[1295][16],mul_out[1295][17],mul_out[1295][18],conv_out[431]);



mul_8x8bit m3888 (image[464],filter[0],mul_out[1296][16]);
mul_8x8bit m3889 (image[465],filter[1],mul_out[1296][17]);
mul_8x8bit m3890 (image[466],filter[2],mul_out[1296][18]);
mul_8x8bit m3891 (image[492],filter[3],mul_out[1297][16]);
mul_8x8bit m3892 (image[493],filter[4],mul_out[1297][17]);
mul_8x8bit m3893 (image[494],filter[5],mul_out[1297][18]);
mul_8x8bit m3894 (image[520],filter[6],mul_out[1298][16]);
mul_8x8bit m3895 (image[521],filter[7],mul_out[1298][17]);
mul_8x8bit m3896 (image[522],filter[8],mul_out[1298][18]);

adder_8bit ad432 (mul_out[1296][16],mul_out[1296][17],mul_out[1296][18],mul_out[1297][16],mul_out[1297][17],mul_out[1297][18],mul_out[1298][16],mul_out[1298][17],mul_out[1298][18],conv_out[432]);



mul_8x8bit m3897 (image[465],filter[0],mul_out[1299][16]);
mul_8x8bit m3898 (image[466],filter[1],mul_out[1299][17]);
mul_8x8bit m3899 (image[467],filter[2],mul_out[1299][18]);
mul_8x8bit m3900 (image[493],filter[3],mul_out[1300][16]);
mul_8x8bit m3901 (image[494],filter[4],mul_out[1300][17]);
mul_8x8bit m3902 (image[495],filter[5],mul_out[1300][18]);
mul_8x8bit m3903 (image[521],filter[6],mul_out[1301][16]);
mul_8x8bit m3904 (image[522],filter[7],mul_out[1301][17]);
mul_8x8bit m3905 (image[523],filter[8],mul_out[1301][18]);

adder_8bit ad433 (mul_out[1299][16],mul_out[1299][17],mul_out[1299][18],mul_out[1300][16],mul_out[1300][17],mul_out[1300][18],mul_out[1301][16],mul_out[1301][17],mul_out[1301][18],conv_out[433]);



mul_8x8bit m3906 (image[466],filter[0],mul_out[1302][16]);
mul_8x8bit m3907 (image[467],filter[1],mul_out[1302][17]);
mul_8x8bit m3908 (image[468],filter[2],mul_out[1302][18]);
mul_8x8bit m3909 (image[494],filter[3],mul_out[1303][16]);
mul_8x8bit m3910 (image[495],filter[4],mul_out[1303][17]);
mul_8x8bit m3911 (image[496],filter[5],mul_out[1303][18]);
mul_8x8bit m3912 (image[522],filter[6],mul_out[1304][16]);
mul_8x8bit m3913 (image[523],filter[7],mul_out[1304][17]);
mul_8x8bit m3914 (image[524],filter[8],mul_out[1304][18]);

adder_8bit ad434 (mul_out[1302][16],mul_out[1302][17],mul_out[1302][18],mul_out[1303][16],mul_out[1303][17],mul_out[1303][18],mul_out[1304][16],mul_out[1304][17],mul_out[1304][18],conv_out[434]);



mul_8x8bit m3915 (image[467],filter[0],mul_out[1305][16]);
mul_8x8bit m3916 (image[468],filter[1],mul_out[1305][17]);
mul_8x8bit m3917 (image[469],filter[2],mul_out[1305][18]);
mul_8x8bit m3918 (image[495],filter[3],mul_out[1306][16]);
mul_8x8bit m3919 (image[496],filter[4],mul_out[1306][17]);
mul_8x8bit m3920 (image[497],filter[5],mul_out[1306][18]);
mul_8x8bit m3921 (image[523],filter[6],mul_out[1307][16]);
mul_8x8bit m3922 (image[524],filter[7],mul_out[1307][17]);
mul_8x8bit m3923 (image[525],filter[8],mul_out[1307][18]);

adder_8bit ad435 (mul_out[1305][16],mul_out[1305][17],mul_out[1305][18],mul_out[1306][16],mul_out[1306][17],mul_out[1306][18],mul_out[1307][16],mul_out[1307][17],mul_out[1307][18],conv_out[435]);



mul_8x8bit m3924 (image[468],filter[0],mul_out[1308][16]);
mul_8x8bit m3925 (image[469],filter[1],mul_out[1308][17]);
mul_8x8bit m3926 (image[470],filter[2],mul_out[1308][18]);
mul_8x8bit m3927 (image[496],filter[3],mul_out[1309][16]);
mul_8x8bit m3928 (image[497],filter[4],mul_out[1309][17]);
mul_8x8bit m3929 (image[498],filter[5],mul_out[1309][18]);
mul_8x8bit m3930 (image[524],filter[6],mul_out[1310][16]);
mul_8x8bit m3931 (image[525],filter[7],mul_out[1310][17]);
mul_8x8bit m3932 (image[526],filter[8],mul_out[1310][18]);

adder_8bit ad436 (mul_out[1308][16],mul_out[1308][17],mul_out[1308][18],mul_out[1309][16],mul_out[1309][17],mul_out[1309][18],mul_out[1310][16],mul_out[1310][17],mul_out[1310][18],conv_out[436]);



mul_8x8bit m3933 (image[469],filter[0],mul_out[1311][16]);
mul_8x8bit m3934 (image[470],filter[1],mul_out[1311][17]);
mul_8x8bit m3935 (image[471],filter[2],mul_out[1311][18]);
mul_8x8bit m3936 (image[497],filter[3],mul_out[1312][16]);
mul_8x8bit m3937 (image[498],filter[4],mul_out[1312][17]);
mul_8x8bit m3938 (image[499],filter[5],mul_out[1312][18]);
mul_8x8bit m3939 (image[525],filter[6],mul_out[1313][16]);
mul_8x8bit m3940 (image[526],filter[7],mul_out[1313][17]);
mul_8x8bit m3941 (image[527],filter[8],mul_out[1313][18]);

adder_8bit ad437 (mul_out[1311][16],mul_out[1311][17],mul_out[1311][18],mul_out[1312][16],mul_out[1312][17],mul_out[1312][18],mul_out[1313][16],mul_out[1313][17],mul_out[1313][18],conv_out[437]);



mul_8x8bit m3942 (image[470],filter[0],mul_out[1314][16]);
mul_8x8bit m3943 (image[471],filter[1],mul_out[1314][17]);
mul_8x8bit m3944 (image[472],filter[2],mul_out[1314][18]);
mul_8x8bit m3945 (image[498],filter[3],mul_out[1315][16]);
mul_8x8bit m3946 (image[499],filter[4],mul_out[1315][17]);
mul_8x8bit m3947 (image[500],filter[5],mul_out[1315][18]);
mul_8x8bit m3948 (image[526],filter[6],mul_out[1316][16]);
mul_8x8bit m3949 (image[527],filter[7],mul_out[1316][17]);
mul_8x8bit m3950 (image[528],filter[8],mul_out[1316][18]);

adder_8bit ad438 (mul_out[1314][16],mul_out[1314][17],mul_out[1314][18],mul_out[1315][16],mul_out[1315][17],mul_out[1315][18],mul_out[1316][16],mul_out[1316][17],mul_out[1316][18],conv_out[438]);



mul_8x8bit m3951 (image[471],filter[0],mul_out[1317][16]);
mul_8x8bit m3952 (image[472],filter[1],mul_out[1317][17]);
mul_8x8bit m3953 (image[473],filter[2],mul_out[1317][18]);
mul_8x8bit m3954 (image[499],filter[3],mul_out[1318][16]);
mul_8x8bit m3955 (image[500],filter[4],mul_out[1318][17]);
mul_8x8bit m3956 (image[501],filter[5],mul_out[1318][18]);
mul_8x8bit m3957 (image[527],filter[6],mul_out[1319][16]);
mul_8x8bit m3958 (image[528],filter[7],mul_out[1319][17]);
mul_8x8bit m3959 (image[529],filter[8],mul_out[1319][18]);

adder_8bit ad439 (mul_out[1317][16],mul_out[1317][17],mul_out[1317][18],mul_out[1318][16],mul_out[1318][17],mul_out[1318][18],mul_out[1319][16],mul_out[1319][17],mul_out[1319][18],conv_out[439]);



mul_8x8bit m3960 (image[472],filter[0],mul_out[1320][16]);
mul_8x8bit m3961 (image[473],filter[1],mul_out[1320][17]);
mul_8x8bit m3962 (image[474],filter[2],mul_out[1320][18]);
mul_8x8bit m3963 (image[500],filter[3],mul_out[1321][16]);
mul_8x8bit m3964 (image[501],filter[4],mul_out[1321][17]);
mul_8x8bit m3965 (image[502],filter[5],mul_out[1321][18]);
mul_8x8bit m3966 (image[528],filter[6],mul_out[1322][16]);
mul_8x8bit m3967 (image[529],filter[7],mul_out[1322][17]);
mul_8x8bit m3968 (image[530],filter[8],mul_out[1322][18]);

adder_8bit ad440 (mul_out[1320][16],mul_out[1320][17],mul_out[1320][18],mul_out[1321][16],mul_out[1321][17],mul_out[1321][18],mul_out[1322][16],mul_out[1322][17],mul_out[1322][18],conv_out[440]);



mul_8x8bit m3969 (image[473],filter[0],mul_out[1323][16]);
mul_8x8bit m3970 (image[474],filter[1],mul_out[1323][17]);
mul_8x8bit m3971 (image[475],filter[2],mul_out[1323][18]);
mul_8x8bit m3972 (image[501],filter[3],mul_out[1324][16]);
mul_8x8bit m3973 (image[502],filter[4],mul_out[1324][17]);
mul_8x8bit m3974 (image[503],filter[5],mul_out[1324][18]);
mul_8x8bit m3975 (image[529],filter[6],mul_out[1325][16]);
mul_8x8bit m3976 (image[530],filter[7],mul_out[1325][17]);
mul_8x8bit m3977 (image[531],filter[8],mul_out[1325][18]);

adder_8bit ad441 (mul_out[1323][16],mul_out[1323][17],mul_out[1323][18],mul_out[1324][16],mul_out[1324][17],mul_out[1324][18],mul_out[1325][16],mul_out[1325][17],mul_out[1325][18],conv_out[441]);



mul_8x8bit m3978 (image[476],filter[0],mul_out[1326][17]);
mul_8x8bit m3979 (image[477],filter[1],mul_out[1326][18]);
mul_8x8bit m3980 (image[478],filter[2],mul_out[1326][19]);
mul_8x8bit m3981 (image[504],filter[3],mul_out[1327][17]);
mul_8x8bit m3982 (image[505],filter[4],mul_out[1327][18]);
mul_8x8bit m3983 (image[506],filter[5],mul_out[1327][19]);
mul_8x8bit m3984 (image[532],filter[6],mul_out[1328][17]);
mul_8x8bit m3985 (image[533],filter[7],mul_out[1328][18]);
mul_8x8bit m3986 (image[534],filter[8],mul_out[1328][19]);

adder_8bit ad442 (mul_out[1326][17],mul_out[1326][18],mul_out[1326][19],mul_out[1327][17],mul_out[1327][18],mul_out[1327][19],mul_out[1328][17],mul_out[1328][18],mul_out[1328][19],conv_out[442]);



mul_8x8bit m3987 (image[477],filter[0],mul_out[1329][17]);
mul_8x8bit m3988 (image[478],filter[1],mul_out[1329][18]);
mul_8x8bit m3989 (image[479],filter[2],mul_out[1329][19]);
mul_8x8bit m3990 (image[505],filter[3],mul_out[1330][17]);
mul_8x8bit m3991 (image[506],filter[4],mul_out[1330][18]);
mul_8x8bit m3992 (image[507],filter[5],mul_out[1330][19]);
mul_8x8bit m3993 (image[533],filter[6],mul_out[1331][17]);
mul_8x8bit m3994 (image[534],filter[7],mul_out[1331][18]);
mul_8x8bit m3995 (image[535],filter[8],mul_out[1331][19]);

adder_8bit ad443 (mul_out[1329][17],mul_out[1329][18],mul_out[1329][19],mul_out[1330][17],mul_out[1330][18],mul_out[1330][19],mul_out[1331][17],mul_out[1331][18],mul_out[1331][19],conv_out[443]);



mul_8x8bit m3996 (image[478],filter[0],mul_out[1332][17]);
mul_8x8bit m3997 (image[479],filter[1],mul_out[1332][18]);
mul_8x8bit m3998 (image[480],filter[2],mul_out[1332][19]);
mul_8x8bit m3999 (image[506],filter[3],mul_out[1333][17]);
mul_8x8bit m4000 (image[507],filter[4],mul_out[1333][18]);
mul_8x8bit m4001 (image[508],filter[5],mul_out[1333][19]);
mul_8x8bit m4002 (image[534],filter[6],mul_out[1334][17]);
mul_8x8bit m4003 (image[535],filter[7],mul_out[1334][18]);
mul_8x8bit m4004 (image[536],filter[8],mul_out[1334][19]);

adder_8bit ad444 (mul_out[1332][17],mul_out[1332][18],mul_out[1332][19],mul_out[1333][17],mul_out[1333][18],mul_out[1333][19],mul_out[1334][17],mul_out[1334][18],mul_out[1334][19],conv_out[444]);



mul_8x8bit m4005 (image[479],filter[0],mul_out[1335][17]);
mul_8x8bit m4006 (image[480],filter[1],mul_out[1335][18]);
mul_8x8bit m4007 (image[481],filter[2],mul_out[1335][19]);
mul_8x8bit m4008 (image[507],filter[3],mul_out[1336][17]);
mul_8x8bit m4009 (image[508],filter[4],mul_out[1336][18]);
mul_8x8bit m4010 (image[509],filter[5],mul_out[1336][19]);
mul_8x8bit m4011 (image[535],filter[6],mul_out[1337][17]);
mul_8x8bit m4012 (image[536],filter[7],mul_out[1337][18]);
mul_8x8bit m4013 (image[537],filter[8],mul_out[1337][19]);

adder_8bit ad445 (mul_out[1335][17],mul_out[1335][18],mul_out[1335][19],mul_out[1336][17],mul_out[1336][18],mul_out[1336][19],mul_out[1337][17],mul_out[1337][18],mul_out[1337][19],conv_out[445]);



mul_8x8bit m4014 (image[480],filter[0],mul_out[1338][17]);
mul_8x8bit m4015 (image[481],filter[1],mul_out[1338][18]);
mul_8x8bit m4016 (image[482],filter[2],mul_out[1338][19]);
mul_8x8bit m4017 (image[508],filter[3],mul_out[1339][17]);
mul_8x8bit m4018 (image[509],filter[4],mul_out[1339][18]);
mul_8x8bit m4019 (image[510],filter[5],mul_out[1339][19]);
mul_8x8bit m4020 (image[536],filter[6],mul_out[1340][17]);
mul_8x8bit m4021 (image[537],filter[7],mul_out[1340][18]);
mul_8x8bit m4022 (image[538],filter[8],mul_out[1340][19]);

adder_8bit ad446 (mul_out[1338][17],mul_out[1338][18],mul_out[1338][19],mul_out[1339][17],mul_out[1339][18],mul_out[1339][19],mul_out[1340][17],mul_out[1340][18],mul_out[1340][19],conv_out[446]);



mul_8x8bit m4023 (image[481],filter[0],mul_out[1341][17]);
mul_8x8bit m4024 (image[482],filter[1],mul_out[1341][18]);
mul_8x8bit m4025 (image[483],filter[2],mul_out[1341][19]);
mul_8x8bit m4026 (image[509],filter[3],mul_out[1342][17]);
mul_8x8bit m4027 (image[510],filter[4],mul_out[1342][18]);
mul_8x8bit m4028 (image[511],filter[5],mul_out[1342][19]);
mul_8x8bit m4029 (image[537],filter[6],mul_out[1343][17]);
mul_8x8bit m4030 (image[538],filter[7],mul_out[1343][18]);
mul_8x8bit m4031 (image[539],filter[8],mul_out[1343][19]);

adder_8bit ad447 (mul_out[1341][17],mul_out[1341][18],mul_out[1341][19],mul_out[1342][17],mul_out[1342][18],mul_out[1342][19],mul_out[1343][17],mul_out[1343][18],mul_out[1343][19],conv_out[447]);



mul_8x8bit m4032 (image[482],filter[0],mul_out[1344][17]);
mul_8x8bit m4033 (image[483],filter[1],mul_out[1344][18]);
mul_8x8bit m4034 (image[484],filter[2],mul_out[1344][19]);
mul_8x8bit m4035 (image[510],filter[3],mul_out[1345][17]);
mul_8x8bit m4036 (image[511],filter[4],mul_out[1345][18]);
mul_8x8bit m4037 (image[512],filter[5],mul_out[1345][19]);
mul_8x8bit m4038 (image[538],filter[6],mul_out[1346][17]);
mul_8x8bit m4039 (image[539],filter[7],mul_out[1346][18]);
mul_8x8bit m4040 (image[540],filter[8],mul_out[1346][19]);

adder_8bit ad448 (mul_out[1344][17],mul_out[1344][18],mul_out[1344][19],mul_out[1345][17],mul_out[1345][18],mul_out[1345][19],mul_out[1346][17],mul_out[1346][18],mul_out[1346][19],conv_out[448]);



mul_8x8bit m4041 (image[483],filter[0],mul_out[1347][17]);
mul_8x8bit m4042 (image[484],filter[1],mul_out[1347][18]);
mul_8x8bit m4043 (image[485],filter[2],mul_out[1347][19]);
mul_8x8bit m4044 (image[511],filter[3],mul_out[1348][17]);
mul_8x8bit m4045 (image[512],filter[4],mul_out[1348][18]);
mul_8x8bit m4046 (image[513],filter[5],mul_out[1348][19]);
mul_8x8bit m4047 (image[539],filter[6],mul_out[1349][17]);
mul_8x8bit m4048 (image[540],filter[7],mul_out[1349][18]);
mul_8x8bit m4049 (image[541],filter[8],mul_out[1349][19]);

adder_8bit ad449 (mul_out[1347][17],mul_out[1347][18],mul_out[1347][19],mul_out[1348][17],mul_out[1348][18],mul_out[1348][19],mul_out[1349][17],mul_out[1349][18],mul_out[1349][19],conv_out[449]);



mul_8x8bit m4050 (image[484],filter[0],mul_out[1350][17]);
mul_8x8bit m4051 (image[485],filter[1],mul_out[1350][18]);
mul_8x8bit m4052 (image[486],filter[2],mul_out[1350][19]);
mul_8x8bit m4053 (image[512],filter[3],mul_out[1351][17]);
mul_8x8bit m4054 (image[513],filter[4],mul_out[1351][18]);
mul_8x8bit m4055 (image[514],filter[5],mul_out[1351][19]);
mul_8x8bit m4056 (image[540],filter[6],mul_out[1352][17]);
mul_8x8bit m4057 (image[541],filter[7],mul_out[1352][18]);
mul_8x8bit m4058 (image[542],filter[8],mul_out[1352][19]);

adder_8bit ad450 (mul_out[1350][17],mul_out[1350][18],mul_out[1350][19],mul_out[1351][17],mul_out[1351][18],mul_out[1351][19],mul_out[1352][17],mul_out[1352][18],mul_out[1352][19],conv_out[450]);



mul_8x8bit m4059 (image[485],filter[0],mul_out[1353][17]);
mul_8x8bit m4060 (image[486],filter[1],mul_out[1353][18]);
mul_8x8bit m4061 (image[487],filter[2],mul_out[1353][19]);
mul_8x8bit m4062 (image[513],filter[3],mul_out[1354][17]);
mul_8x8bit m4063 (image[514],filter[4],mul_out[1354][18]);
mul_8x8bit m4064 (image[515],filter[5],mul_out[1354][19]);
mul_8x8bit m4065 (image[541],filter[6],mul_out[1355][17]);
mul_8x8bit m4066 (image[542],filter[7],mul_out[1355][18]);
mul_8x8bit m4067 (image[543],filter[8],mul_out[1355][19]);

adder_8bit ad451 (mul_out[1353][17],mul_out[1353][18],mul_out[1353][19],mul_out[1354][17],mul_out[1354][18],mul_out[1354][19],mul_out[1355][17],mul_out[1355][18],mul_out[1355][19],conv_out[451]);



mul_8x8bit m4068 (image[486],filter[0],mul_out[1356][17]);
mul_8x8bit m4069 (image[487],filter[1],mul_out[1356][18]);
mul_8x8bit m4070 (image[488],filter[2],mul_out[1356][19]);
mul_8x8bit m4071 (image[514],filter[3],mul_out[1357][17]);
mul_8x8bit m4072 (image[515],filter[4],mul_out[1357][18]);
mul_8x8bit m4073 (image[516],filter[5],mul_out[1357][19]);
mul_8x8bit m4074 (image[542],filter[6],mul_out[1358][17]);
mul_8x8bit m4075 (image[543],filter[7],mul_out[1358][18]);
mul_8x8bit m4076 (image[544],filter[8],mul_out[1358][19]);

adder_8bit ad452 (mul_out[1356][17],mul_out[1356][18],mul_out[1356][19],mul_out[1357][17],mul_out[1357][18],mul_out[1357][19],mul_out[1358][17],mul_out[1358][18],mul_out[1358][19],conv_out[452]);



mul_8x8bit m4077 (image[487],filter[0],mul_out[1359][17]);
mul_8x8bit m4078 (image[488],filter[1],mul_out[1359][18]);
mul_8x8bit m4079 (image[489],filter[2],mul_out[1359][19]);
mul_8x8bit m4080 (image[515],filter[3],mul_out[1360][17]);
mul_8x8bit m4081 (image[516],filter[4],mul_out[1360][18]);
mul_8x8bit m4082 (image[517],filter[5],mul_out[1360][19]);
mul_8x8bit m4083 (image[543],filter[6],mul_out[1361][17]);
mul_8x8bit m4084 (image[544],filter[7],mul_out[1361][18]);
mul_8x8bit m4085 (image[545],filter[8],mul_out[1361][19]);

adder_8bit ad453 (mul_out[1359][17],mul_out[1359][18],mul_out[1359][19],mul_out[1360][17],mul_out[1360][18],mul_out[1360][19],mul_out[1361][17],mul_out[1361][18],mul_out[1361][19],conv_out[453]);



mul_8x8bit m4086 (image[488],filter[0],mul_out[1362][17]);
mul_8x8bit m4087 (image[489],filter[1],mul_out[1362][18]);
mul_8x8bit m4088 (image[490],filter[2],mul_out[1362][19]);
mul_8x8bit m4089 (image[516],filter[3],mul_out[1363][17]);
mul_8x8bit m4090 (image[517],filter[4],mul_out[1363][18]);
mul_8x8bit m4091 (image[518],filter[5],mul_out[1363][19]);
mul_8x8bit m4092 (image[544],filter[6],mul_out[1364][17]);
mul_8x8bit m4093 (image[545],filter[7],mul_out[1364][18]);
mul_8x8bit m4094 (image[546],filter[8],mul_out[1364][19]);

adder_8bit ad454 (mul_out[1362][17],mul_out[1362][18],mul_out[1362][19],mul_out[1363][17],mul_out[1363][18],mul_out[1363][19],mul_out[1364][17],mul_out[1364][18],mul_out[1364][19],conv_out[454]);



mul_8x8bit m4095 (image[489],filter[0],mul_out[1365][17]);
mul_8x8bit m4096 (image[490],filter[1],mul_out[1365][18]);
mul_8x8bit m4097 (image[491],filter[2],mul_out[1365][19]);
mul_8x8bit m4098 (image[517],filter[3],mul_out[1366][17]);
mul_8x8bit m4099 (image[518],filter[4],mul_out[1366][18]);
mul_8x8bit m4100 (image[519],filter[5],mul_out[1366][19]);
mul_8x8bit m4101 (image[545],filter[6],mul_out[1367][17]);
mul_8x8bit m4102 (image[546],filter[7],mul_out[1367][18]);
mul_8x8bit m4103 (image[547],filter[8],mul_out[1367][19]);

adder_8bit ad455 (mul_out[1365][17],mul_out[1365][18],mul_out[1365][19],mul_out[1366][17],mul_out[1366][18],mul_out[1366][19],mul_out[1367][17],mul_out[1367][18],mul_out[1367][19],conv_out[455]);



mul_8x8bit m4104 (image[490],filter[0],mul_out[1368][17]);
mul_8x8bit m4105 (image[491],filter[1],mul_out[1368][18]);
mul_8x8bit m4106 (image[492],filter[2],mul_out[1368][19]);
mul_8x8bit m4107 (image[518],filter[3],mul_out[1369][17]);
mul_8x8bit m4108 (image[519],filter[4],mul_out[1369][18]);
mul_8x8bit m4109 (image[520],filter[5],mul_out[1369][19]);
mul_8x8bit m4110 (image[546],filter[6],mul_out[1370][17]);
mul_8x8bit m4111 (image[547],filter[7],mul_out[1370][18]);
mul_8x8bit m4112 (image[548],filter[8],mul_out[1370][19]);

adder_8bit ad456 (mul_out[1368][17],mul_out[1368][18],mul_out[1368][19],mul_out[1369][17],mul_out[1369][18],mul_out[1369][19],mul_out[1370][17],mul_out[1370][18],mul_out[1370][19],conv_out[456]);



mul_8x8bit m4113 (image[491],filter[0],mul_out[1371][17]);
mul_8x8bit m4114 (image[492],filter[1],mul_out[1371][18]);
mul_8x8bit m4115 (image[493],filter[2],mul_out[1371][19]);
mul_8x8bit m4116 (image[519],filter[3],mul_out[1372][17]);
mul_8x8bit m4117 (image[520],filter[4],mul_out[1372][18]);
mul_8x8bit m4118 (image[521],filter[5],mul_out[1372][19]);
mul_8x8bit m4119 (image[547],filter[6],mul_out[1373][17]);
mul_8x8bit m4120 (image[548],filter[7],mul_out[1373][18]);
mul_8x8bit m4121 (image[549],filter[8],mul_out[1373][19]);

adder_8bit ad457 (mul_out[1371][17],mul_out[1371][18],mul_out[1371][19],mul_out[1372][17],mul_out[1372][18],mul_out[1372][19],mul_out[1373][17],mul_out[1373][18],mul_out[1373][19],conv_out[457]);



mul_8x8bit m4122 (image[492],filter[0],mul_out[1374][17]);
mul_8x8bit m4123 (image[493],filter[1],mul_out[1374][18]);
mul_8x8bit m4124 (image[494],filter[2],mul_out[1374][19]);
mul_8x8bit m4125 (image[520],filter[3],mul_out[1375][17]);
mul_8x8bit m4126 (image[521],filter[4],mul_out[1375][18]);
mul_8x8bit m4127 (image[522],filter[5],mul_out[1375][19]);
mul_8x8bit m4128 (image[548],filter[6],mul_out[1376][17]);
mul_8x8bit m4129 (image[549],filter[7],mul_out[1376][18]);
mul_8x8bit m4130 (image[550],filter[8],mul_out[1376][19]);

adder_8bit ad458 (mul_out[1374][17],mul_out[1374][18],mul_out[1374][19],mul_out[1375][17],mul_out[1375][18],mul_out[1375][19],mul_out[1376][17],mul_out[1376][18],mul_out[1376][19],conv_out[458]);



mul_8x8bit m4131 (image[493],filter[0],mul_out[1377][17]);
mul_8x8bit m4132 (image[494],filter[1],mul_out[1377][18]);
mul_8x8bit m4133 (image[495],filter[2],mul_out[1377][19]);
mul_8x8bit m4134 (image[521],filter[3],mul_out[1378][17]);
mul_8x8bit m4135 (image[522],filter[4],mul_out[1378][18]);
mul_8x8bit m4136 (image[523],filter[5],mul_out[1378][19]);
mul_8x8bit m4137 (image[549],filter[6],mul_out[1379][17]);
mul_8x8bit m4138 (image[550],filter[7],mul_out[1379][18]);
mul_8x8bit m4139 (image[551],filter[8],mul_out[1379][19]);

adder_8bit ad459 (mul_out[1377][17],mul_out[1377][18],mul_out[1377][19],mul_out[1378][17],mul_out[1378][18],mul_out[1378][19],mul_out[1379][17],mul_out[1379][18],mul_out[1379][19],conv_out[459]);



mul_8x8bit m4140 (image[494],filter[0],mul_out[1380][17]);
mul_8x8bit m4141 (image[495],filter[1],mul_out[1380][18]);
mul_8x8bit m4142 (image[496],filter[2],mul_out[1380][19]);
mul_8x8bit m4143 (image[522],filter[3],mul_out[1381][17]);
mul_8x8bit m4144 (image[523],filter[4],mul_out[1381][18]);
mul_8x8bit m4145 (image[524],filter[5],mul_out[1381][19]);
mul_8x8bit m4146 (image[550],filter[6],mul_out[1382][17]);
mul_8x8bit m4147 (image[551],filter[7],mul_out[1382][18]);
mul_8x8bit m4148 (image[552],filter[8],mul_out[1382][19]);

adder_8bit ad460 (mul_out[1380][17],mul_out[1380][18],mul_out[1380][19],mul_out[1381][17],mul_out[1381][18],mul_out[1381][19],mul_out[1382][17],mul_out[1382][18],mul_out[1382][19],conv_out[460]);



mul_8x8bit m4149 (image[495],filter[0],mul_out[1383][17]);
mul_8x8bit m4150 (image[496],filter[1],mul_out[1383][18]);
mul_8x8bit m4151 (image[497],filter[2],mul_out[1383][19]);
mul_8x8bit m4152 (image[523],filter[3],mul_out[1384][17]);
mul_8x8bit m4153 (image[524],filter[4],mul_out[1384][18]);
mul_8x8bit m4154 (image[525],filter[5],mul_out[1384][19]);
mul_8x8bit m4155 (image[551],filter[6],mul_out[1385][17]);
mul_8x8bit m4156 (image[552],filter[7],mul_out[1385][18]);
mul_8x8bit m4157 (image[553],filter[8],mul_out[1385][19]);

adder_8bit ad461 (mul_out[1383][17],mul_out[1383][18],mul_out[1383][19],mul_out[1384][17],mul_out[1384][18],mul_out[1384][19],mul_out[1385][17],mul_out[1385][18],mul_out[1385][19],conv_out[461]);



mul_8x8bit m4158 (image[496],filter[0],mul_out[1386][17]);
mul_8x8bit m4159 (image[497],filter[1],mul_out[1386][18]);
mul_8x8bit m4160 (image[498],filter[2],mul_out[1386][19]);
mul_8x8bit m4161 (image[524],filter[3],mul_out[1387][17]);
mul_8x8bit m4162 (image[525],filter[4],mul_out[1387][18]);
mul_8x8bit m4163 (image[526],filter[5],mul_out[1387][19]);
mul_8x8bit m4164 (image[552],filter[6],mul_out[1388][17]);
mul_8x8bit m4165 (image[553],filter[7],mul_out[1388][18]);
mul_8x8bit m4166 (image[554],filter[8],mul_out[1388][19]);

adder_8bit ad462 (mul_out[1386][17],mul_out[1386][18],mul_out[1386][19],mul_out[1387][17],mul_out[1387][18],mul_out[1387][19],mul_out[1388][17],mul_out[1388][18],mul_out[1388][19],conv_out[462]);



mul_8x8bit m4167 (image[497],filter[0],mul_out[1389][17]);
mul_8x8bit m4168 (image[498],filter[1],mul_out[1389][18]);
mul_8x8bit m4169 (image[499],filter[2],mul_out[1389][19]);
mul_8x8bit m4170 (image[525],filter[3],mul_out[1390][17]);
mul_8x8bit m4171 (image[526],filter[4],mul_out[1390][18]);
mul_8x8bit m4172 (image[527],filter[5],mul_out[1390][19]);
mul_8x8bit m4173 (image[553],filter[6],mul_out[1391][17]);
mul_8x8bit m4174 (image[554],filter[7],mul_out[1391][18]);
mul_8x8bit m4175 (image[555],filter[8],mul_out[1391][19]);

adder_8bit ad463 (mul_out[1389][17],mul_out[1389][18],mul_out[1389][19],mul_out[1390][17],mul_out[1390][18],mul_out[1390][19],mul_out[1391][17],mul_out[1391][18],mul_out[1391][19],conv_out[463]);



mul_8x8bit m4176 (image[498],filter[0],mul_out[1392][17]);
mul_8x8bit m4177 (image[499],filter[1],mul_out[1392][18]);
mul_8x8bit m4178 (image[500],filter[2],mul_out[1392][19]);
mul_8x8bit m4179 (image[526],filter[3],mul_out[1393][17]);
mul_8x8bit m4180 (image[527],filter[4],mul_out[1393][18]);
mul_8x8bit m4181 (image[528],filter[5],mul_out[1393][19]);
mul_8x8bit m4182 (image[554],filter[6],mul_out[1394][17]);
mul_8x8bit m4183 (image[555],filter[7],mul_out[1394][18]);
mul_8x8bit m4184 (image[556],filter[8],mul_out[1394][19]);

adder_8bit ad464 (mul_out[1392][17],mul_out[1392][18],mul_out[1392][19],mul_out[1393][17],mul_out[1393][18],mul_out[1393][19],mul_out[1394][17],mul_out[1394][18],mul_out[1394][19],conv_out[464]);



mul_8x8bit m4185 (image[499],filter[0],mul_out[1395][17]);
mul_8x8bit m4186 (image[500],filter[1],mul_out[1395][18]);
mul_8x8bit m4187 (image[501],filter[2],mul_out[1395][19]);
mul_8x8bit m4188 (image[527],filter[3],mul_out[1396][17]);
mul_8x8bit m4189 (image[528],filter[4],mul_out[1396][18]);
mul_8x8bit m4190 (image[529],filter[5],mul_out[1396][19]);
mul_8x8bit m4191 (image[555],filter[6],mul_out[1397][17]);
mul_8x8bit m4192 (image[556],filter[7],mul_out[1397][18]);
mul_8x8bit m4193 (image[557],filter[8],mul_out[1397][19]);

adder_8bit ad465 (mul_out[1395][17],mul_out[1395][18],mul_out[1395][19],mul_out[1396][17],mul_out[1396][18],mul_out[1396][19],mul_out[1397][17],mul_out[1397][18],mul_out[1397][19],conv_out[465]);



mul_8x8bit m4194 (image[500],filter[0],mul_out[1398][17]);
mul_8x8bit m4195 (image[501],filter[1],mul_out[1398][18]);
mul_8x8bit m4196 (image[502],filter[2],mul_out[1398][19]);
mul_8x8bit m4197 (image[528],filter[3],mul_out[1399][17]);
mul_8x8bit m4198 (image[529],filter[4],mul_out[1399][18]);
mul_8x8bit m4199 (image[530],filter[5],mul_out[1399][19]);
mul_8x8bit m4200 (image[556],filter[6],mul_out[1400][17]);
mul_8x8bit m4201 (image[557],filter[7],mul_out[1400][18]);
mul_8x8bit m4202 (image[558],filter[8],mul_out[1400][19]);

adder_8bit ad466 (mul_out[1398][17],mul_out[1398][18],mul_out[1398][19],mul_out[1399][17],mul_out[1399][18],mul_out[1399][19],mul_out[1400][17],mul_out[1400][18],mul_out[1400][19],conv_out[466]);



mul_8x8bit m4203 (image[501],filter[0],mul_out[1401][17]);
mul_8x8bit m4204 (image[502],filter[1],mul_out[1401][18]);
mul_8x8bit m4205 (image[503],filter[2],mul_out[1401][19]);
mul_8x8bit m4206 (image[529],filter[3],mul_out[1402][17]);
mul_8x8bit m4207 (image[530],filter[4],mul_out[1402][18]);
mul_8x8bit m4208 (image[531],filter[5],mul_out[1402][19]);
mul_8x8bit m4209 (image[557],filter[6],mul_out[1403][17]);
mul_8x8bit m4210 (image[558],filter[7],mul_out[1403][18]);
mul_8x8bit m4211 (image[559],filter[8],mul_out[1403][19]);

adder_8bit ad467 (mul_out[1401][17],mul_out[1401][18],mul_out[1401][19],mul_out[1402][17],mul_out[1402][18],mul_out[1402][19],mul_out[1403][17],mul_out[1403][18],mul_out[1403][19],conv_out[467]);



mul_8x8bit m4212 (image[504],filter[0],mul_out[1404][18]);
mul_8x8bit m4213 (image[505],filter[1],mul_out[1404][19]);
mul_8x8bit m4214 (image[506],filter[2],mul_out[1404][20]);
mul_8x8bit m4215 (image[532],filter[3],mul_out[1405][18]);
mul_8x8bit m4216 (image[533],filter[4],mul_out[1405][19]);
mul_8x8bit m4217 (image[534],filter[5],mul_out[1405][20]);
mul_8x8bit m4218 (image[560],filter[6],mul_out[1406][18]);
mul_8x8bit m4219 (image[561],filter[7],mul_out[1406][19]);
mul_8x8bit m4220 (image[562],filter[8],mul_out[1406][20]);

adder_8bit ad468 (mul_out[1404][18],mul_out[1404][19],mul_out[1404][20],mul_out[1405][18],mul_out[1405][19],mul_out[1405][20],mul_out[1406][18],mul_out[1406][19],mul_out[1406][20],conv_out[468]);



mul_8x8bit m4221 (image[505],filter[0],mul_out[1407][18]);
mul_8x8bit m4222 (image[506],filter[1],mul_out[1407][19]);
mul_8x8bit m4223 (image[507],filter[2],mul_out[1407][20]);
mul_8x8bit m4224 (image[533],filter[3],mul_out[1408][18]);
mul_8x8bit m4225 (image[534],filter[4],mul_out[1408][19]);
mul_8x8bit m4226 (image[535],filter[5],mul_out[1408][20]);
mul_8x8bit m4227 (image[561],filter[6],mul_out[1409][18]);
mul_8x8bit m4228 (image[562],filter[7],mul_out[1409][19]);
mul_8x8bit m4229 (image[563],filter[8],mul_out[1409][20]);

adder_8bit ad469 (mul_out[1407][18],mul_out[1407][19],mul_out[1407][20],mul_out[1408][18],mul_out[1408][19],mul_out[1408][20],mul_out[1409][18],mul_out[1409][19],mul_out[1409][20],conv_out[469]);



mul_8x8bit m4230 (image[506],filter[0],mul_out[1410][18]);
mul_8x8bit m4231 (image[507],filter[1],mul_out[1410][19]);
mul_8x8bit m4232 (image[508],filter[2],mul_out[1410][20]);
mul_8x8bit m4233 (image[534],filter[3],mul_out[1411][18]);
mul_8x8bit m4234 (image[535],filter[4],mul_out[1411][19]);
mul_8x8bit m4235 (image[536],filter[5],mul_out[1411][20]);
mul_8x8bit m4236 (image[562],filter[6],mul_out[1412][18]);
mul_8x8bit m4237 (image[563],filter[7],mul_out[1412][19]);
mul_8x8bit m4238 (image[564],filter[8],mul_out[1412][20]);

adder_8bit ad470 (mul_out[1410][18],mul_out[1410][19],mul_out[1410][20],mul_out[1411][18],mul_out[1411][19],mul_out[1411][20],mul_out[1412][18],mul_out[1412][19],mul_out[1412][20],conv_out[470]);



mul_8x8bit m4239 (image[507],filter[0],mul_out[1413][18]);
mul_8x8bit m4240 (image[508],filter[1],mul_out[1413][19]);
mul_8x8bit m4241 (image[509],filter[2],mul_out[1413][20]);
mul_8x8bit m4242 (image[535],filter[3],mul_out[1414][18]);
mul_8x8bit m4243 (image[536],filter[4],mul_out[1414][19]);
mul_8x8bit m4244 (image[537],filter[5],mul_out[1414][20]);
mul_8x8bit m4245 (image[563],filter[6],mul_out[1415][18]);
mul_8x8bit m4246 (image[564],filter[7],mul_out[1415][19]);
mul_8x8bit m4247 (image[565],filter[8],mul_out[1415][20]);

adder_8bit ad471 (mul_out[1413][18],mul_out[1413][19],mul_out[1413][20],mul_out[1414][18],mul_out[1414][19],mul_out[1414][20],mul_out[1415][18],mul_out[1415][19],mul_out[1415][20],conv_out[471]);



mul_8x8bit m4248 (image[508],filter[0],mul_out[1416][18]);
mul_8x8bit m4249 (image[509],filter[1],mul_out[1416][19]);
mul_8x8bit m4250 (image[510],filter[2],mul_out[1416][20]);
mul_8x8bit m4251 (image[536],filter[3],mul_out[1417][18]);
mul_8x8bit m4252 (image[537],filter[4],mul_out[1417][19]);
mul_8x8bit m4253 (image[538],filter[5],mul_out[1417][20]);
mul_8x8bit m4254 (image[564],filter[6],mul_out[1418][18]);
mul_8x8bit m4255 (image[565],filter[7],mul_out[1418][19]);
mul_8x8bit m4256 (image[566],filter[8],mul_out[1418][20]);

adder_8bit ad472 (mul_out[1416][18],mul_out[1416][19],mul_out[1416][20],mul_out[1417][18],mul_out[1417][19],mul_out[1417][20],mul_out[1418][18],mul_out[1418][19],mul_out[1418][20],conv_out[472]);



mul_8x8bit m4257 (image[509],filter[0],mul_out[1419][18]);
mul_8x8bit m4258 (image[510],filter[1],mul_out[1419][19]);
mul_8x8bit m4259 (image[511],filter[2],mul_out[1419][20]);
mul_8x8bit m4260 (image[537],filter[3],mul_out[1420][18]);
mul_8x8bit m4261 (image[538],filter[4],mul_out[1420][19]);
mul_8x8bit m4262 (image[539],filter[5],mul_out[1420][20]);
mul_8x8bit m4263 (image[565],filter[6],mul_out[1421][18]);
mul_8x8bit m4264 (image[566],filter[7],mul_out[1421][19]);
mul_8x8bit m4265 (image[567],filter[8],mul_out[1421][20]);

adder_8bit ad473 (mul_out[1419][18],mul_out[1419][19],mul_out[1419][20],mul_out[1420][18],mul_out[1420][19],mul_out[1420][20],mul_out[1421][18],mul_out[1421][19],mul_out[1421][20],conv_out[473]);



mul_8x8bit m4266 (image[510],filter[0],mul_out[1422][18]);
mul_8x8bit m4267 (image[511],filter[1],mul_out[1422][19]);
mul_8x8bit m4268 (image[512],filter[2],mul_out[1422][20]);
mul_8x8bit m4269 (image[538],filter[3],mul_out[1423][18]);
mul_8x8bit m4270 (image[539],filter[4],mul_out[1423][19]);
mul_8x8bit m4271 (image[540],filter[5],mul_out[1423][20]);
mul_8x8bit m4272 (image[566],filter[6],mul_out[1424][18]);
mul_8x8bit m4273 (image[567],filter[7],mul_out[1424][19]);
mul_8x8bit m4274 (image[568],filter[8],mul_out[1424][20]);

adder_8bit ad474 (mul_out[1422][18],mul_out[1422][19],mul_out[1422][20],mul_out[1423][18],mul_out[1423][19],mul_out[1423][20],mul_out[1424][18],mul_out[1424][19],mul_out[1424][20],conv_out[474]);



mul_8x8bit m4275 (image[511],filter[0],mul_out[1425][18]);
mul_8x8bit m4276 (image[512],filter[1],mul_out[1425][19]);
mul_8x8bit m4277 (image[513],filter[2],mul_out[1425][20]);
mul_8x8bit m4278 (image[539],filter[3],mul_out[1426][18]);
mul_8x8bit m4279 (image[540],filter[4],mul_out[1426][19]);
mul_8x8bit m4280 (image[541],filter[5],mul_out[1426][20]);
mul_8x8bit m4281 (image[567],filter[6],mul_out[1427][18]);
mul_8x8bit m4282 (image[568],filter[7],mul_out[1427][19]);
mul_8x8bit m4283 (image[569],filter[8],mul_out[1427][20]);

adder_8bit ad475 (mul_out[1425][18],mul_out[1425][19],mul_out[1425][20],mul_out[1426][18],mul_out[1426][19],mul_out[1426][20],mul_out[1427][18],mul_out[1427][19],mul_out[1427][20],conv_out[475]);



mul_8x8bit m4284 (image[512],filter[0],mul_out[1428][18]);
mul_8x8bit m4285 (image[513],filter[1],mul_out[1428][19]);
mul_8x8bit m4286 (image[514],filter[2],mul_out[1428][20]);
mul_8x8bit m4287 (image[540],filter[3],mul_out[1429][18]);
mul_8x8bit m4288 (image[541],filter[4],mul_out[1429][19]);
mul_8x8bit m4289 (image[542],filter[5],mul_out[1429][20]);
mul_8x8bit m4290 (image[568],filter[6],mul_out[1430][18]);
mul_8x8bit m4291 (image[569],filter[7],mul_out[1430][19]);
mul_8x8bit m4292 (image[570],filter[8],mul_out[1430][20]);

adder_8bit ad476 (mul_out[1428][18],mul_out[1428][19],mul_out[1428][20],mul_out[1429][18],mul_out[1429][19],mul_out[1429][20],mul_out[1430][18],mul_out[1430][19],mul_out[1430][20],conv_out[476]);



mul_8x8bit m4293 (image[513],filter[0],mul_out[1431][18]);
mul_8x8bit m4294 (image[514],filter[1],mul_out[1431][19]);
mul_8x8bit m4295 (image[515],filter[2],mul_out[1431][20]);
mul_8x8bit m4296 (image[541],filter[3],mul_out[1432][18]);
mul_8x8bit m4297 (image[542],filter[4],mul_out[1432][19]);
mul_8x8bit m4298 (image[543],filter[5],mul_out[1432][20]);
mul_8x8bit m4299 (image[569],filter[6],mul_out[1433][18]);
mul_8x8bit m4300 (image[570],filter[7],mul_out[1433][19]);
mul_8x8bit m4301 (image[571],filter[8],mul_out[1433][20]);

adder_8bit ad477 (mul_out[1431][18],mul_out[1431][19],mul_out[1431][20],mul_out[1432][18],mul_out[1432][19],mul_out[1432][20],mul_out[1433][18],mul_out[1433][19],mul_out[1433][20],conv_out[477]);



mul_8x8bit m4302 (image[514],filter[0],mul_out[1434][18]);
mul_8x8bit m4303 (image[515],filter[1],mul_out[1434][19]);
mul_8x8bit m4304 (image[516],filter[2],mul_out[1434][20]);
mul_8x8bit m4305 (image[542],filter[3],mul_out[1435][18]);
mul_8x8bit m4306 (image[543],filter[4],mul_out[1435][19]);
mul_8x8bit m4307 (image[544],filter[5],mul_out[1435][20]);
mul_8x8bit m4308 (image[570],filter[6],mul_out[1436][18]);
mul_8x8bit m4309 (image[571],filter[7],mul_out[1436][19]);
mul_8x8bit m4310 (image[572],filter[8],mul_out[1436][20]);

adder_8bit ad478 (mul_out[1434][18],mul_out[1434][19],mul_out[1434][20],mul_out[1435][18],mul_out[1435][19],mul_out[1435][20],mul_out[1436][18],mul_out[1436][19],mul_out[1436][20],conv_out[478]);



mul_8x8bit m4311 (image[515],filter[0],mul_out[1437][18]);
mul_8x8bit m4312 (image[516],filter[1],mul_out[1437][19]);
mul_8x8bit m4313 (image[517],filter[2],mul_out[1437][20]);
mul_8x8bit m4314 (image[543],filter[3],mul_out[1438][18]);
mul_8x8bit m4315 (image[544],filter[4],mul_out[1438][19]);
mul_8x8bit m4316 (image[545],filter[5],mul_out[1438][20]);
mul_8x8bit m4317 (image[571],filter[6],mul_out[1439][18]);
mul_8x8bit m4318 (image[572],filter[7],mul_out[1439][19]);
mul_8x8bit m4319 (image[573],filter[8],mul_out[1439][20]);

adder_8bit ad479 (mul_out[1437][18],mul_out[1437][19],mul_out[1437][20],mul_out[1438][18],mul_out[1438][19],mul_out[1438][20],mul_out[1439][18],mul_out[1439][19],mul_out[1439][20],conv_out[479]);



mul_8x8bit m4320 (image[516],filter[0],mul_out[1440][18]);
mul_8x8bit m4321 (image[517],filter[1],mul_out[1440][19]);
mul_8x8bit m4322 (image[518],filter[2],mul_out[1440][20]);
mul_8x8bit m4323 (image[544],filter[3],mul_out[1441][18]);
mul_8x8bit m4324 (image[545],filter[4],mul_out[1441][19]);
mul_8x8bit m4325 (image[546],filter[5],mul_out[1441][20]);
mul_8x8bit m4326 (image[572],filter[6],mul_out[1442][18]);
mul_8x8bit m4327 (image[573],filter[7],mul_out[1442][19]);
mul_8x8bit m4328 (image[574],filter[8],mul_out[1442][20]);

adder_8bit ad480 (mul_out[1440][18],mul_out[1440][19],mul_out[1440][20],mul_out[1441][18],mul_out[1441][19],mul_out[1441][20],mul_out[1442][18],mul_out[1442][19],mul_out[1442][20],conv_out[480]);



mul_8x8bit m4329 (image[517],filter[0],mul_out[1443][18]);
mul_8x8bit m4330 (image[518],filter[1],mul_out[1443][19]);
mul_8x8bit m4331 (image[519],filter[2],mul_out[1443][20]);
mul_8x8bit m4332 (image[545],filter[3],mul_out[1444][18]);
mul_8x8bit m4333 (image[546],filter[4],mul_out[1444][19]);
mul_8x8bit m4334 (image[547],filter[5],mul_out[1444][20]);
mul_8x8bit m4335 (image[573],filter[6],mul_out[1445][18]);
mul_8x8bit m4336 (image[574],filter[7],mul_out[1445][19]);
mul_8x8bit m4337 (image[575],filter[8],mul_out[1445][20]);

adder_8bit ad481 (mul_out[1443][18],mul_out[1443][19],mul_out[1443][20],mul_out[1444][18],mul_out[1444][19],mul_out[1444][20],mul_out[1445][18],mul_out[1445][19],mul_out[1445][20],conv_out[481]);



mul_8x8bit m4338 (image[518],filter[0],mul_out[1446][18]);
mul_8x8bit m4339 (image[519],filter[1],mul_out[1446][19]);
mul_8x8bit m4340 (image[520],filter[2],mul_out[1446][20]);
mul_8x8bit m4341 (image[546],filter[3],mul_out[1447][18]);
mul_8x8bit m4342 (image[547],filter[4],mul_out[1447][19]);
mul_8x8bit m4343 (image[548],filter[5],mul_out[1447][20]);
mul_8x8bit m4344 (image[574],filter[6],mul_out[1448][18]);
mul_8x8bit m4345 (image[575],filter[7],mul_out[1448][19]);
mul_8x8bit m4346 (image[576],filter[8],mul_out[1448][20]);

adder_8bit ad482 (mul_out[1446][18],mul_out[1446][19],mul_out[1446][20],mul_out[1447][18],mul_out[1447][19],mul_out[1447][20],mul_out[1448][18],mul_out[1448][19],mul_out[1448][20],conv_out[482]);



mul_8x8bit m4347 (image[519],filter[0],mul_out[1449][18]);
mul_8x8bit m4348 (image[520],filter[1],mul_out[1449][19]);
mul_8x8bit m4349 (image[521],filter[2],mul_out[1449][20]);
mul_8x8bit m4350 (image[547],filter[3],mul_out[1450][18]);
mul_8x8bit m4351 (image[548],filter[4],mul_out[1450][19]);
mul_8x8bit m4352 (image[549],filter[5],mul_out[1450][20]);
mul_8x8bit m4353 (image[575],filter[6],mul_out[1451][18]);
mul_8x8bit m4354 (image[576],filter[7],mul_out[1451][19]);
mul_8x8bit m4355 (image[577],filter[8],mul_out[1451][20]);

adder_8bit ad483 (mul_out[1449][18],mul_out[1449][19],mul_out[1449][20],mul_out[1450][18],mul_out[1450][19],mul_out[1450][20],mul_out[1451][18],mul_out[1451][19],mul_out[1451][20],conv_out[483]);



mul_8x8bit m4356 (image[520],filter[0],mul_out[1452][18]);
mul_8x8bit m4357 (image[521],filter[1],mul_out[1452][19]);
mul_8x8bit m4358 (image[522],filter[2],mul_out[1452][20]);
mul_8x8bit m4359 (image[548],filter[3],mul_out[1453][18]);
mul_8x8bit m4360 (image[549],filter[4],mul_out[1453][19]);
mul_8x8bit m4361 (image[550],filter[5],mul_out[1453][20]);
mul_8x8bit m4362 (image[576],filter[6],mul_out[1454][18]);
mul_8x8bit m4363 (image[577],filter[7],mul_out[1454][19]);
mul_8x8bit m4364 (image[578],filter[8],mul_out[1454][20]);

adder_8bit ad484 (mul_out[1452][18],mul_out[1452][19],mul_out[1452][20],mul_out[1453][18],mul_out[1453][19],mul_out[1453][20],mul_out[1454][18],mul_out[1454][19],mul_out[1454][20],conv_out[484]);



mul_8x8bit m4365 (image[521],filter[0],mul_out[1455][18]);
mul_8x8bit m4366 (image[522],filter[1],mul_out[1455][19]);
mul_8x8bit m4367 (image[523],filter[2],mul_out[1455][20]);
mul_8x8bit m4368 (image[549],filter[3],mul_out[1456][18]);
mul_8x8bit m4369 (image[550],filter[4],mul_out[1456][19]);
mul_8x8bit m4370 (image[551],filter[5],mul_out[1456][20]);
mul_8x8bit m4371 (image[577],filter[6],mul_out[1457][18]);
mul_8x8bit m4372 (image[578],filter[7],mul_out[1457][19]);
mul_8x8bit m4373 (image[579],filter[8],mul_out[1457][20]);

adder_8bit ad485 (mul_out[1455][18],mul_out[1455][19],mul_out[1455][20],mul_out[1456][18],mul_out[1456][19],mul_out[1456][20],mul_out[1457][18],mul_out[1457][19],mul_out[1457][20],conv_out[485]);



mul_8x8bit m4374 (image[522],filter[0],mul_out[1458][18]);
mul_8x8bit m4375 (image[523],filter[1],mul_out[1458][19]);
mul_8x8bit m4376 (image[524],filter[2],mul_out[1458][20]);
mul_8x8bit m4377 (image[550],filter[3],mul_out[1459][18]);
mul_8x8bit m4378 (image[551],filter[4],mul_out[1459][19]);
mul_8x8bit m4379 (image[552],filter[5],mul_out[1459][20]);
mul_8x8bit m4380 (image[578],filter[6],mul_out[1460][18]);
mul_8x8bit m4381 (image[579],filter[7],mul_out[1460][19]);
mul_8x8bit m4382 (image[580],filter[8],mul_out[1460][20]);

adder_8bit ad486 (mul_out[1458][18],mul_out[1458][19],mul_out[1458][20],mul_out[1459][18],mul_out[1459][19],mul_out[1459][20],mul_out[1460][18],mul_out[1460][19],mul_out[1460][20],conv_out[486]);



mul_8x8bit m4383 (image[523],filter[0],mul_out[1461][18]);
mul_8x8bit m4384 (image[524],filter[1],mul_out[1461][19]);
mul_8x8bit m4385 (image[525],filter[2],mul_out[1461][20]);
mul_8x8bit m4386 (image[551],filter[3],mul_out[1462][18]);
mul_8x8bit m4387 (image[552],filter[4],mul_out[1462][19]);
mul_8x8bit m4388 (image[553],filter[5],mul_out[1462][20]);
mul_8x8bit m4389 (image[579],filter[6],mul_out[1463][18]);
mul_8x8bit m4390 (image[580],filter[7],mul_out[1463][19]);
mul_8x8bit m4391 (image[581],filter[8],mul_out[1463][20]);

adder_8bit ad487 (mul_out[1461][18],mul_out[1461][19],mul_out[1461][20],mul_out[1462][18],mul_out[1462][19],mul_out[1462][20],mul_out[1463][18],mul_out[1463][19],mul_out[1463][20],conv_out[487]);



mul_8x8bit m4392 (image[524],filter[0],mul_out[1464][18]);
mul_8x8bit m4393 (image[525],filter[1],mul_out[1464][19]);
mul_8x8bit m4394 (image[526],filter[2],mul_out[1464][20]);
mul_8x8bit m4395 (image[552],filter[3],mul_out[1465][18]);
mul_8x8bit m4396 (image[553],filter[4],mul_out[1465][19]);
mul_8x8bit m4397 (image[554],filter[5],mul_out[1465][20]);
mul_8x8bit m4398 (image[580],filter[6],mul_out[1466][18]);
mul_8x8bit m4399 (image[581],filter[7],mul_out[1466][19]);
mul_8x8bit m4400 (image[582],filter[8],mul_out[1466][20]);

adder_8bit ad488 (mul_out[1464][18],mul_out[1464][19],mul_out[1464][20],mul_out[1465][18],mul_out[1465][19],mul_out[1465][20],mul_out[1466][18],mul_out[1466][19],mul_out[1466][20],conv_out[488]);



mul_8x8bit m4401 (image[525],filter[0],mul_out[1467][18]);
mul_8x8bit m4402 (image[526],filter[1],mul_out[1467][19]);
mul_8x8bit m4403 (image[527],filter[2],mul_out[1467][20]);
mul_8x8bit m4404 (image[553],filter[3],mul_out[1468][18]);
mul_8x8bit m4405 (image[554],filter[4],mul_out[1468][19]);
mul_8x8bit m4406 (image[555],filter[5],mul_out[1468][20]);
mul_8x8bit m4407 (image[581],filter[6],mul_out[1469][18]);
mul_8x8bit m4408 (image[582],filter[7],mul_out[1469][19]);
mul_8x8bit m4409 (image[583],filter[8],mul_out[1469][20]);

adder_8bit ad489 (mul_out[1467][18],mul_out[1467][19],mul_out[1467][20],mul_out[1468][18],mul_out[1468][19],mul_out[1468][20],mul_out[1469][18],mul_out[1469][19],mul_out[1469][20],conv_out[489]);



mul_8x8bit m4410 (image[526],filter[0],mul_out[1470][18]);
mul_8x8bit m4411 (image[527],filter[1],mul_out[1470][19]);
mul_8x8bit m4412 (image[528],filter[2],mul_out[1470][20]);
mul_8x8bit m4413 (image[554],filter[3],mul_out[1471][18]);
mul_8x8bit m4414 (image[555],filter[4],mul_out[1471][19]);
mul_8x8bit m4415 (image[556],filter[5],mul_out[1471][20]);
mul_8x8bit m4416 (image[582],filter[6],mul_out[1472][18]);
mul_8x8bit m4417 (image[583],filter[7],mul_out[1472][19]);
mul_8x8bit m4418 (image[584],filter[8],mul_out[1472][20]);

adder_8bit ad490 (mul_out[1470][18],mul_out[1470][19],mul_out[1470][20],mul_out[1471][18],mul_out[1471][19],mul_out[1471][20],mul_out[1472][18],mul_out[1472][19],mul_out[1472][20],conv_out[490]);



mul_8x8bit m4419 (image[527],filter[0],mul_out[1473][18]);
mul_8x8bit m4420 (image[528],filter[1],mul_out[1473][19]);
mul_8x8bit m4421 (image[529],filter[2],mul_out[1473][20]);
mul_8x8bit m4422 (image[555],filter[3],mul_out[1474][18]);
mul_8x8bit m4423 (image[556],filter[4],mul_out[1474][19]);
mul_8x8bit m4424 (image[557],filter[5],mul_out[1474][20]);
mul_8x8bit m4425 (image[583],filter[6],mul_out[1475][18]);
mul_8x8bit m4426 (image[584],filter[7],mul_out[1475][19]);
mul_8x8bit m4427 (image[585],filter[8],mul_out[1475][20]);

adder_8bit ad491 (mul_out[1473][18],mul_out[1473][19],mul_out[1473][20],mul_out[1474][18],mul_out[1474][19],mul_out[1474][20],mul_out[1475][18],mul_out[1475][19],mul_out[1475][20],conv_out[491]);



mul_8x8bit m4428 (image[528],filter[0],mul_out[1476][18]);
mul_8x8bit m4429 (image[529],filter[1],mul_out[1476][19]);
mul_8x8bit m4430 (image[530],filter[2],mul_out[1476][20]);
mul_8x8bit m4431 (image[556],filter[3],mul_out[1477][18]);
mul_8x8bit m4432 (image[557],filter[4],mul_out[1477][19]);
mul_8x8bit m4433 (image[558],filter[5],mul_out[1477][20]);
mul_8x8bit m4434 (image[584],filter[6],mul_out[1478][18]);
mul_8x8bit m4435 (image[585],filter[7],mul_out[1478][19]);
mul_8x8bit m4436 (image[586],filter[8],mul_out[1478][20]);

adder_8bit ad492 (mul_out[1476][18],mul_out[1476][19],mul_out[1476][20],mul_out[1477][18],mul_out[1477][19],mul_out[1477][20],mul_out[1478][18],mul_out[1478][19],mul_out[1478][20],conv_out[492]);



mul_8x8bit m4437 (image[529],filter[0],mul_out[1479][18]);
mul_8x8bit m4438 (image[530],filter[1],mul_out[1479][19]);
mul_8x8bit m4439 (image[531],filter[2],mul_out[1479][20]);
mul_8x8bit m4440 (image[557],filter[3],mul_out[1480][18]);
mul_8x8bit m4441 (image[558],filter[4],mul_out[1480][19]);
mul_8x8bit m4442 (image[559],filter[5],mul_out[1480][20]);
mul_8x8bit m4443 (image[585],filter[6],mul_out[1481][18]);
mul_8x8bit m4444 (image[586],filter[7],mul_out[1481][19]);
mul_8x8bit m4445 (image[587],filter[8],mul_out[1481][20]);

adder_8bit ad493 (mul_out[1479][18],mul_out[1479][19],mul_out[1479][20],mul_out[1480][18],mul_out[1480][19],mul_out[1480][20],mul_out[1481][18],mul_out[1481][19],mul_out[1481][20],conv_out[493]);



mul_8x8bit m4446 (image[532],filter[0],mul_out[1482][19]);
mul_8x8bit m4447 (image[533],filter[1],mul_out[1482][20]);
mul_8x8bit m4448 (image[534],filter[2],mul_out[1482][21]);
mul_8x8bit m4449 (image[560],filter[3],mul_out[1483][19]);
mul_8x8bit m4450 (image[561],filter[4],mul_out[1483][20]);
mul_8x8bit m4451 (image[562],filter[5],mul_out[1483][21]);
mul_8x8bit m4452 (image[588],filter[6],mul_out[1484][19]);
mul_8x8bit m4453 (image[589],filter[7],mul_out[1484][20]);
mul_8x8bit m4454 (image[590],filter[8],mul_out[1484][21]);

adder_8bit ad494 (mul_out[1482][19],mul_out[1482][20],mul_out[1482][21],mul_out[1483][19],mul_out[1483][20],mul_out[1483][21],mul_out[1484][19],mul_out[1484][20],mul_out[1484][21],conv_out[494]);



mul_8x8bit m4455 (image[533],filter[0],mul_out[1485][19]);
mul_8x8bit m4456 (image[534],filter[1],mul_out[1485][20]);
mul_8x8bit m4457 (image[535],filter[2],mul_out[1485][21]);
mul_8x8bit m4458 (image[561],filter[3],mul_out[1486][19]);
mul_8x8bit m4459 (image[562],filter[4],mul_out[1486][20]);
mul_8x8bit m4460 (image[563],filter[5],mul_out[1486][21]);
mul_8x8bit m4461 (image[589],filter[6],mul_out[1487][19]);
mul_8x8bit m4462 (image[590],filter[7],mul_out[1487][20]);
mul_8x8bit m4463 (image[591],filter[8],mul_out[1487][21]);

adder_8bit ad495 (mul_out[1485][19],mul_out[1485][20],mul_out[1485][21],mul_out[1486][19],mul_out[1486][20],mul_out[1486][21],mul_out[1487][19],mul_out[1487][20],mul_out[1487][21],conv_out[495]);



mul_8x8bit m4464 (image[534],filter[0],mul_out[1488][19]);
mul_8x8bit m4465 (image[535],filter[1],mul_out[1488][20]);
mul_8x8bit m4466 (image[536],filter[2],mul_out[1488][21]);
mul_8x8bit m4467 (image[562],filter[3],mul_out[1489][19]);
mul_8x8bit m4468 (image[563],filter[4],mul_out[1489][20]);
mul_8x8bit m4469 (image[564],filter[5],mul_out[1489][21]);
mul_8x8bit m4470 (image[590],filter[6],mul_out[1490][19]);
mul_8x8bit m4471 (image[591],filter[7],mul_out[1490][20]);
mul_8x8bit m4472 (image[592],filter[8],mul_out[1490][21]);

adder_8bit ad496 (mul_out[1488][19],mul_out[1488][20],mul_out[1488][21],mul_out[1489][19],mul_out[1489][20],mul_out[1489][21],mul_out[1490][19],mul_out[1490][20],mul_out[1490][21],conv_out[496]);



mul_8x8bit m4473 (image[535],filter[0],mul_out[1491][19]);
mul_8x8bit m4474 (image[536],filter[1],mul_out[1491][20]);
mul_8x8bit m4475 (image[537],filter[2],mul_out[1491][21]);
mul_8x8bit m4476 (image[563],filter[3],mul_out[1492][19]);
mul_8x8bit m4477 (image[564],filter[4],mul_out[1492][20]);
mul_8x8bit m4478 (image[565],filter[5],mul_out[1492][21]);
mul_8x8bit m4479 (image[591],filter[6],mul_out[1493][19]);
mul_8x8bit m4480 (image[592],filter[7],mul_out[1493][20]);
mul_8x8bit m4481 (image[593],filter[8],mul_out[1493][21]);

adder_8bit ad497 (mul_out[1491][19],mul_out[1491][20],mul_out[1491][21],mul_out[1492][19],mul_out[1492][20],mul_out[1492][21],mul_out[1493][19],mul_out[1493][20],mul_out[1493][21],conv_out[497]);



mul_8x8bit m4482 (image[536],filter[0],mul_out[1494][19]);
mul_8x8bit m4483 (image[537],filter[1],mul_out[1494][20]);
mul_8x8bit m4484 (image[538],filter[2],mul_out[1494][21]);
mul_8x8bit m4485 (image[564],filter[3],mul_out[1495][19]);
mul_8x8bit m4486 (image[565],filter[4],mul_out[1495][20]);
mul_8x8bit m4487 (image[566],filter[5],mul_out[1495][21]);
mul_8x8bit m4488 (image[592],filter[6],mul_out[1496][19]);
mul_8x8bit m4489 (image[593],filter[7],mul_out[1496][20]);
mul_8x8bit m4490 (image[594],filter[8],mul_out[1496][21]);

adder_8bit ad498 (mul_out[1494][19],mul_out[1494][20],mul_out[1494][21],mul_out[1495][19],mul_out[1495][20],mul_out[1495][21],mul_out[1496][19],mul_out[1496][20],mul_out[1496][21],conv_out[498]);



mul_8x8bit m4491 (image[537],filter[0],mul_out[1497][19]);
mul_8x8bit m4492 (image[538],filter[1],mul_out[1497][20]);
mul_8x8bit m4493 (image[539],filter[2],mul_out[1497][21]);
mul_8x8bit m4494 (image[565],filter[3],mul_out[1498][19]);
mul_8x8bit m4495 (image[566],filter[4],mul_out[1498][20]);
mul_8x8bit m4496 (image[567],filter[5],mul_out[1498][21]);
mul_8x8bit m4497 (image[593],filter[6],mul_out[1499][19]);
mul_8x8bit m4498 (image[594],filter[7],mul_out[1499][20]);
mul_8x8bit m4499 (image[595],filter[8],mul_out[1499][21]);

adder_8bit ad499 (mul_out[1497][19],mul_out[1497][20],mul_out[1497][21],mul_out[1498][19],mul_out[1498][20],mul_out[1498][21],mul_out[1499][19],mul_out[1499][20],mul_out[1499][21],conv_out[499]);



mul_8x8bit m4500 (image[538],filter[0],mul_out[1500][19]);
mul_8x8bit m4501 (image[539],filter[1],mul_out[1500][20]);
mul_8x8bit m4502 (image[540],filter[2],mul_out[1500][21]);
mul_8x8bit m4503 (image[566],filter[3],mul_out[1501][19]);
mul_8x8bit m4504 (image[567],filter[4],mul_out[1501][20]);
mul_8x8bit m4505 (image[568],filter[5],mul_out[1501][21]);
mul_8x8bit m4506 (image[594],filter[6],mul_out[1502][19]);
mul_8x8bit m4507 (image[595],filter[7],mul_out[1502][20]);
mul_8x8bit m4508 (image[596],filter[8],mul_out[1502][21]);

adder_8bit ad500 (mul_out[1500][19],mul_out[1500][20],mul_out[1500][21],mul_out[1501][19],mul_out[1501][20],mul_out[1501][21],mul_out[1502][19],mul_out[1502][20],mul_out[1502][21],conv_out[500]);



mul_8x8bit m4509 (image[539],filter[0],mul_out[1503][19]);
mul_8x8bit m4510 (image[540],filter[1],mul_out[1503][20]);
mul_8x8bit m4511 (image[541],filter[2],mul_out[1503][21]);
mul_8x8bit m4512 (image[567],filter[3],mul_out[1504][19]);
mul_8x8bit m4513 (image[568],filter[4],mul_out[1504][20]);
mul_8x8bit m4514 (image[569],filter[5],mul_out[1504][21]);
mul_8x8bit m4515 (image[595],filter[6],mul_out[1505][19]);
mul_8x8bit m4516 (image[596],filter[7],mul_out[1505][20]);
mul_8x8bit m4517 (image[597],filter[8],mul_out[1505][21]);

adder_8bit ad501 (mul_out[1503][19],mul_out[1503][20],mul_out[1503][21],mul_out[1504][19],mul_out[1504][20],mul_out[1504][21],mul_out[1505][19],mul_out[1505][20],mul_out[1505][21],conv_out[501]);



mul_8x8bit m4518 (image[540],filter[0],mul_out[1506][19]);
mul_8x8bit m4519 (image[541],filter[1],mul_out[1506][20]);
mul_8x8bit m4520 (image[542],filter[2],mul_out[1506][21]);
mul_8x8bit m4521 (image[568],filter[3],mul_out[1507][19]);
mul_8x8bit m4522 (image[569],filter[4],mul_out[1507][20]);
mul_8x8bit m4523 (image[570],filter[5],mul_out[1507][21]);
mul_8x8bit m4524 (image[596],filter[6],mul_out[1508][19]);
mul_8x8bit m4525 (image[597],filter[7],mul_out[1508][20]);
mul_8x8bit m4526 (image[598],filter[8],mul_out[1508][21]);

adder_8bit ad502 (mul_out[1506][19],mul_out[1506][20],mul_out[1506][21],mul_out[1507][19],mul_out[1507][20],mul_out[1507][21],mul_out[1508][19],mul_out[1508][20],mul_out[1508][21],conv_out[502]);



mul_8x8bit m4527 (image[541],filter[0],mul_out[1509][19]);
mul_8x8bit m4528 (image[542],filter[1],mul_out[1509][20]);
mul_8x8bit m4529 (image[543],filter[2],mul_out[1509][21]);
mul_8x8bit m4530 (image[569],filter[3],mul_out[1510][19]);
mul_8x8bit m4531 (image[570],filter[4],mul_out[1510][20]);
mul_8x8bit m4532 (image[571],filter[5],mul_out[1510][21]);
mul_8x8bit m4533 (image[597],filter[6],mul_out[1511][19]);
mul_8x8bit m4534 (image[598],filter[7],mul_out[1511][20]);
mul_8x8bit m4535 (image[599],filter[8],mul_out[1511][21]);

adder_8bit ad503 (mul_out[1509][19],mul_out[1509][20],mul_out[1509][21],mul_out[1510][19],mul_out[1510][20],mul_out[1510][21],mul_out[1511][19],mul_out[1511][20],mul_out[1511][21],conv_out[503]);



mul_8x8bit m4536 (image[542],filter[0],mul_out[1512][19]);
mul_8x8bit m4537 (image[543],filter[1],mul_out[1512][20]);
mul_8x8bit m4538 (image[544],filter[2],mul_out[1512][21]);
mul_8x8bit m4539 (image[570],filter[3],mul_out[1513][19]);
mul_8x8bit m4540 (image[571],filter[4],mul_out[1513][20]);
mul_8x8bit m4541 (image[572],filter[5],mul_out[1513][21]);
mul_8x8bit m4542 (image[598],filter[6],mul_out[1514][19]);
mul_8x8bit m4543 (image[599],filter[7],mul_out[1514][20]);
mul_8x8bit m4544 (image[600],filter[8],mul_out[1514][21]);

adder_8bit ad504 (mul_out[1512][19],mul_out[1512][20],mul_out[1512][21],mul_out[1513][19],mul_out[1513][20],mul_out[1513][21],mul_out[1514][19],mul_out[1514][20],mul_out[1514][21],conv_out[504]);



mul_8x8bit m4545 (image[543],filter[0],mul_out[1515][19]);
mul_8x8bit m4546 (image[544],filter[1],mul_out[1515][20]);
mul_8x8bit m4547 (image[545],filter[2],mul_out[1515][21]);
mul_8x8bit m4548 (image[571],filter[3],mul_out[1516][19]);
mul_8x8bit m4549 (image[572],filter[4],mul_out[1516][20]);
mul_8x8bit m4550 (image[573],filter[5],mul_out[1516][21]);
mul_8x8bit m4551 (image[599],filter[6],mul_out[1517][19]);
mul_8x8bit m4552 (image[600],filter[7],mul_out[1517][20]);
mul_8x8bit m4553 (image[601],filter[8],mul_out[1517][21]);

adder_8bit ad505 (mul_out[1515][19],mul_out[1515][20],mul_out[1515][21],mul_out[1516][19],mul_out[1516][20],mul_out[1516][21],mul_out[1517][19],mul_out[1517][20],mul_out[1517][21],conv_out[505]);



mul_8x8bit m4554 (image[544],filter[0],mul_out[1518][19]);
mul_8x8bit m4555 (image[545],filter[1],mul_out[1518][20]);
mul_8x8bit m4556 (image[546],filter[2],mul_out[1518][21]);
mul_8x8bit m4557 (image[572],filter[3],mul_out[1519][19]);
mul_8x8bit m4558 (image[573],filter[4],mul_out[1519][20]);
mul_8x8bit m4559 (image[574],filter[5],mul_out[1519][21]);
mul_8x8bit m4560 (image[600],filter[6],mul_out[1520][19]);
mul_8x8bit m4561 (image[601],filter[7],mul_out[1520][20]);
mul_8x8bit m4562 (image[602],filter[8],mul_out[1520][21]);

adder_8bit ad506 (mul_out[1518][19],mul_out[1518][20],mul_out[1518][21],mul_out[1519][19],mul_out[1519][20],mul_out[1519][21],mul_out[1520][19],mul_out[1520][20],mul_out[1520][21],conv_out[506]);



mul_8x8bit m4563 (image[545],filter[0],mul_out[1521][19]);
mul_8x8bit m4564 (image[546],filter[1],mul_out[1521][20]);
mul_8x8bit m4565 (image[547],filter[2],mul_out[1521][21]);
mul_8x8bit m4566 (image[573],filter[3],mul_out[1522][19]);
mul_8x8bit m4567 (image[574],filter[4],mul_out[1522][20]);
mul_8x8bit m4568 (image[575],filter[5],mul_out[1522][21]);
mul_8x8bit m4569 (image[601],filter[6],mul_out[1523][19]);
mul_8x8bit m4570 (image[602],filter[7],mul_out[1523][20]);
mul_8x8bit m4571 (image[603],filter[8],mul_out[1523][21]);

adder_8bit ad507 (mul_out[1521][19],mul_out[1521][20],mul_out[1521][21],mul_out[1522][19],mul_out[1522][20],mul_out[1522][21],mul_out[1523][19],mul_out[1523][20],mul_out[1523][21],conv_out[507]);



mul_8x8bit m4572 (image[546],filter[0],mul_out[1524][19]);
mul_8x8bit m4573 (image[547],filter[1],mul_out[1524][20]);
mul_8x8bit m4574 (image[548],filter[2],mul_out[1524][21]);
mul_8x8bit m4575 (image[574],filter[3],mul_out[1525][19]);
mul_8x8bit m4576 (image[575],filter[4],mul_out[1525][20]);
mul_8x8bit m4577 (image[576],filter[5],mul_out[1525][21]);
mul_8x8bit m4578 (image[602],filter[6],mul_out[1526][19]);
mul_8x8bit m4579 (image[603],filter[7],mul_out[1526][20]);
mul_8x8bit m4580 (image[604],filter[8],mul_out[1526][21]);

adder_8bit ad508 (mul_out[1524][19],mul_out[1524][20],mul_out[1524][21],mul_out[1525][19],mul_out[1525][20],mul_out[1525][21],mul_out[1526][19],mul_out[1526][20],mul_out[1526][21],conv_out[508]);



mul_8x8bit m4581 (image[547],filter[0],mul_out[1527][19]);
mul_8x8bit m4582 (image[548],filter[1],mul_out[1527][20]);
mul_8x8bit m4583 (image[549],filter[2],mul_out[1527][21]);
mul_8x8bit m4584 (image[575],filter[3],mul_out[1528][19]);
mul_8x8bit m4585 (image[576],filter[4],mul_out[1528][20]);
mul_8x8bit m4586 (image[577],filter[5],mul_out[1528][21]);
mul_8x8bit m4587 (image[603],filter[6],mul_out[1529][19]);
mul_8x8bit m4588 (image[604],filter[7],mul_out[1529][20]);
mul_8x8bit m4589 (image[605],filter[8],mul_out[1529][21]);

adder_8bit ad509 (mul_out[1527][19],mul_out[1527][20],mul_out[1527][21],mul_out[1528][19],mul_out[1528][20],mul_out[1528][21],mul_out[1529][19],mul_out[1529][20],mul_out[1529][21],conv_out[509]);



mul_8x8bit m4590 (image[548],filter[0],mul_out[1530][19]);
mul_8x8bit m4591 (image[549],filter[1],mul_out[1530][20]);
mul_8x8bit m4592 (image[550],filter[2],mul_out[1530][21]);
mul_8x8bit m4593 (image[576],filter[3],mul_out[1531][19]);
mul_8x8bit m4594 (image[577],filter[4],mul_out[1531][20]);
mul_8x8bit m4595 (image[578],filter[5],mul_out[1531][21]);
mul_8x8bit m4596 (image[604],filter[6],mul_out[1532][19]);
mul_8x8bit m4597 (image[605],filter[7],mul_out[1532][20]);
mul_8x8bit m4598 (image[606],filter[8],mul_out[1532][21]);

adder_8bit ad510 (mul_out[1530][19],mul_out[1530][20],mul_out[1530][21],mul_out[1531][19],mul_out[1531][20],mul_out[1531][21],mul_out[1532][19],mul_out[1532][20],mul_out[1532][21],conv_out[510]);



mul_8x8bit m4599 (image[549],filter[0],mul_out[1533][19]);
mul_8x8bit m4600 (image[550],filter[1],mul_out[1533][20]);
mul_8x8bit m4601 (image[551],filter[2],mul_out[1533][21]);
mul_8x8bit m4602 (image[577],filter[3],mul_out[1534][19]);
mul_8x8bit m4603 (image[578],filter[4],mul_out[1534][20]);
mul_8x8bit m4604 (image[579],filter[5],mul_out[1534][21]);
mul_8x8bit m4605 (image[605],filter[6],mul_out[1535][19]);
mul_8x8bit m4606 (image[606],filter[7],mul_out[1535][20]);
mul_8x8bit m4607 (image[607],filter[8],mul_out[1535][21]);

adder_8bit ad511 (mul_out[1533][19],mul_out[1533][20],mul_out[1533][21],mul_out[1534][19],mul_out[1534][20],mul_out[1534][21],mul_out[1535][19],mul_out[1535][20],mul_out[1535][21],conv_out[511]);



mul_8x8bit m4608 (image[550],filter[0],mul_out[1536][19]);
mul_8x8bit m4609 (image[551],filter[1],mul_out[1536][20]);
mul_8x8bit m4610 (image[552],filter[2],mul_out[1536][21]);
mul_8x8bit m4611 (image[578],filter[3],mul_out[1537][19]);
mul_8x8bit m4612 (image[579],filter[4],mul_out[1537][20]);
mul_8x8bit m4613 (image[580],filter[5],mul_out[1537][21]);
mul_8x8bit m4614 (image[606],filter[6],mul_out[1538][19]);
mul_8x8bit m4615 (image[607],filter[7],mul_out[1538][20]);
mul_8x8bit m4616 (image[608],filter[8],mul_out[1538][21]);

adder_8bit ad512 (mul_out[1536][19],mul_out[1536][20],mul_out[1536][21],mul_out[1537][19],mul_out[1537][20],mul_out[1537][21],mul_out[1538][19],mul_out[1538][20],mul_out[1538][21],conv_out[512]);



mul_8x8bit m4617 (image[551],filter[0],mul_out[1539][19]);
mul_8x8bit m4618 (image[552],filter[1],mul_out[1539][20]);
mul_8x8bit m4619 (image[553],filter[2],mul_out[1539][21]);
mul_8x8bit m4620 (image[579],filter[3],mul_out[1540][19]);
mul_8x8bit m4621 (image[580],filter[4],mul_out[1540][20]);
mul_8x8bit m4622 (image[581],filter[5],mul_out[1540][21]);
mul_8x8bit m4623 (image[607],filter[6],mul_out[1541][19]);
mul_8x8bit m4624 (image[608],filter[7],mul_out[1541][20]);
mul_8x8bit m4625 (image[609],filter[8],mul_out[1541][21]);

adder_8bit ad513 (mul_out[1539][19],mul_out[1539][20],mul_out[1539][21],mul_out[1540][19],mul_out[1540][20],mul_out[1540][21],mul_out[1541][19],mul_out[1541][20],mul_out[1541][21],conv_out[513]);



mul_8x8bit m4626 (image[552],filter[0],mul_out[1542][19]);
mul_8x8bit m4627 (image[553],filter[1],mul_out[1542][20]);
mul_8x8bit m4628 (image[554],filter[2],mul_out[1542][21]);
mul_8x8bit m4629 (image[580],filter[3],mul_out[1543][19]);
mul_8x8bit m4630 (image[581],filter[4],mul_out[1543][20]);
mul_8x8bit m4631 (image[582],filter[5],mul_out[1543][21]);
mul_8x8bit m4632 (image[608],filter[6],mul_out[1544][19]);
mul_8x8bit m4633 (image[609],filter[7],mul_out[1544][20]);
mul_8x8bit m4634 (image[610],filter[8],mul_out[1544][21]);

adder_8bit ad514 (mul_out[1542][19],mul_out[1542][20],mul_out[1542][21],mul_out[1543][19],mul_out[1543][20],mul_out[1543][21],mul_out[1544][19],mul_out[1544][20],mul_out[1544][21],conv_out[514]);



mul_8x8bit m4635 (image[553],filter[0],mul_out[1545][19]);
mul_8x8bit m4636 (image[554],filter[1],mul_out[1545][20]);
mul_8x8bit m4637 (image[555],filter[2],mul_out[1545][21]);
mul_8x8bit m4638 (image[581],filter[3],mul_out[1546][19]);
mul_8x8bit m4639 (image[582],filter[4],mul_out[1546][20]);
mul_8x8bit m4640 (image[583],filter[5],mul_out[1546][21]);
mul_8x8bit m4641 (image[609],filter[6],mul_out[1547][19]);
mul_8x8bit m4642 (image[610],filter[7],mul_out[1547][20]);
mul_8x8bit m4643 (image[611],filter[8],mul_out[1547][21]);

adder_8bit ad515 (mul_out[1545][19],mul_out[1545][20],mul_out[1545][21],mul_out[1546][19],mul_out[1546][20],mul_out[1546][21],mul_out[1547][19],mul_out[1547][20],mul_out[1547][21],conv_out[515]);



mul_8x8bit m4644 (image[554],filter[0],mul_out[1548][19]);
mul_8x8bit m4645 (image[555],filter[1],mul_out[1548][20]);
mul_8x8bit m4646 (image[556],filter[2],mul_out[1548][21]);
mul_8x8bit m4647 (image[582],filter[3],mul_out[1549][19]);
mul_8x8bit m4648 (image[583],filter[4],mul_out[1549][20]);
mul_8x8bit m4649 (image[584],filter[5],mul_out[1549][21]);
mul_8x8bit m4650 (image[610],filter[6],mul_out[1550][19]);
mul_8x8bit m4651 (image[611],filter[7],mul_out[1550][20]);
mul_8x8bit m4652 (image[612],filter[8],mul_out[1550][21]);

adder_8bit ad516 (mul_out[1548][19],mul_out[1548][20],mul_out[1548][21],mul_out[1549][19],mul_out[1549][20],mul_out[1549][21],mul_out[1550][19],mul_out[1550][20],mul_out[1550][21],conv_out[516]);



mul_8x8bit m4653 (image[555],filter[0],mul_out[1551][19]);
mul_8x8bit m4654 (image[556],filter[1],mul_out[1551][20]);
mul_8x8bit m4655 (image[557],filter[2],mul_out[1551][21]);
mul_8x8bit m4656 (image[583],filter[3],mul_out[1552][19]);
mul_8x8bit m4657 (image[584],filter[4],mul_out[1552][20]);
mul_8x8bit m4658 (image[585],filter[5],mul_out[1552][21]);
mul_8x8bit m4659 (image[611],filter[6],mul_out[1553][19]);
mul_8x8bit m4660 (image[612],filter[7],mul_out[1553][20]);
mul_8x8bit m4661 (image[613],filter[8],mul_out[1553][21]);

adder_8bit ad517 (mul_out[1551][19],mul_out[1551][20],mul_out[1551][21],mul_out[1552][19],mul_out[1552][20],mul_out[1552][21],mul_out[1553][19],mul_out[1553][20],mul_out[1553][21],conv_out[517]);



mul_8x8bit m4662 (image[556],filter[0],mul_out[1554][19]);
mul_8x8bit m4663 (image[557],filter[1],mul_out[1554][20]);
mul_8x8bit m4664 (image[558],filter[2],mul_out[1554][21]);
mul_8x8bit m4665 (image[584],filter[3],mul_out[1555][19]);
mul_8x8bit m4666 (image[585],filter[4],mul_out[1555][20]);
mul_8x8bit m4667 (image[586],filter[5],mul_out[1555][21]);
mul_8x8bit m4668 (image[612],filter[6],mul_out[1556][19]);
mul_8x8bit m4669 (image[613],filter[7],mul_out[1556][20]);
mul_8x8bit m4670 (image[614],filter[8],mul_out[1556][21]);

adder_8bit ad518 (mul_out[1554][19],mul_out[1554][20],mul_out[1554][21],mul_out[1555][19],mul_out[1555][20],mul_out[1555][21],mul_out[1556][19],mul_out[1556][20],mul_out[1556][21],conv_out[518]);



mul_8x8bit m4671 (image[557],filter[0],mul_out[1557][19]);
mul_8x8bit m4672 (image[558],filter[1],mul_out[1557][20]);
mul_8x8bit m4673 (image[559],filter[2],mul_out[1557][21]);
mul_8x8bit m4674 (image[585],filter[3],mul_out[1558][19]);
mul_8x8bit m4675 (image[586],filter[4],mul_out[1558][20]);
mul_8x8bit m4676 (image[587],filter[5],mul_out[1558][21]);
mul_8x8bit m4677 (image[613],filter[6],mul_out[1559][19]);
mul_8x8bit m4678 (image[614],filter[7],mul_out[1559][20]);
mul_8x8bit m4679 (image[615],filter[8],mul_out[1559][21]);

adder_8bit ad519 (mul_out[1557][19],mul_out[1557][20],mul_out[1557][21],mul_out[1558][19],mul_out[1558][20],mul_out[1558][21],mul_out[1559][19],mul_out[1559][20],mul_out[1559][21],conv_out[519]);



mul_8x8bit m4680 (image[560],filter[0],mul_out[1560][20]);
mul_8x8bit m4681 (image[561],filter[1],mul_out[1560][21]);
mul_8x8bit m4682 (image[562],filter[2],mul_out[1560][22]);
mul_8x8bit m4683 (image[588],filter[3],mul_out[1561][20]);
mul_8x8bit m4684 (image[589],filter[4],mul_out[1561][21]);
mul_8x8bit m4685 (image[590],filter[5],mul_out[1561][22]);
mul_8x8bit m4686 (image[616],filter[6],mul_out[1562][20]);
mul_8x8bit m4687 (image[617],filter[7],mul_out[1562][21]);
mul_8x8bit m4688 (image[618],filter[8],mul_out[1562][22]);

adder_8bit ad520 (mul_out[1560][20],mul_out[1560][21],mul_out[1560][22],mul_out[1561][20],mul_out[1561][21],mul_out[1561][22],mul_out[1562][20],mul_out[1562][21],mul_out[1562][22],conv_out[520]);



mul_8x8bit m4689 (image[561],filter[0],mul_out[1563][20]);
mul_8x8bit m4690 (image[562],filter[1],mul_out[1563][21]);
mul_8x8bit m4691 (image[563],filter[2],mul_out[1563][22]);
mul_8x8bit m4692 (image[589],filter[3],mul_out[1564][20]);
mul_8x8bit m4693 (image[590],filter[4],mul_out[1564][21]);
mul_8x8bit m4694 (image[591],filter[5],mul_out[1564][22]);
mul_8x8bit m4695 (image[617],filter[6],mul_out[1565][20]);
mul_8x8bit m4696 (image[618],filter[7],mul_out[1565][21]);
mul_8x8bit m4697 (image[619],filter[8],mul_out[1565][22]);

adder_8bit ad521 (mul_out[1563][20],mul_out[1563][21],mul_out[1563][22],mul_out[1564][20],mul_out[1564][21],mul_out[1564][22],mul_out[1565][20],mul_out[1565][21],mul_out[1565][22],conv_out[521]);



mul_8x8bit m4698 (image[562],filter[0],mul_out[1566][20]);
mul_8x8bit m4699 (image[563],filter[1],mul_out[1566][21]);
mul_8x8bit m4700 (image[564],filter[2],mul_out[1566][22]);
mul_8x8bit m4701 (image[590],filter[3],mul_out[1567][20]);
mul_8x8bit m4702 (image[591],filter[4],mul_out[1567][21]);
mul_8x8bit m4703 (image[592],filter[5],mul_out[1567][22]);
mul_8x8bit m4704 (image[618],filter[6],mul_out[1568][20]);
mul_8x8bit m4705 (image[619],filter[7],mul_out[1568][21]);
mul_8x8bit m4706 (image[620],filter[8],mul_out[1568][22]);

adder_8bit ad522 (mul_out[1566][20],mul_out[1566][21],mul_out[1566][22],mul_out[1567][20],mul_out[1567][21],mul_out[1567][22],mul_out[1568][20],mul_out[1568][21],mul_out[1568][22],conv_out[522]);



mul_8x8bit m4707 (image[563],filter[0],mul_out[1569][20]);
mul_8x8bit m4708 (image[564],filter[1],mul_out[1569][21]);
mul_8x8bit m4709 (image[565],filter[2],mul_out[1569][22]);
mul_8x8bit m4710 (image[591],filter[3],mul_out[1570][20]);
mul_8x8bit m4711 (image[592],filter[4],mul_out[1570][21]);
mul_8x8bit m4712 (image[593],filter[5],mul_out[1570][22]);
mul_8x8bit m4713 (image[619],filter[6],mul_out[1571][20]);
mul_8x8bit m4714 (image[620],filter[7],mul_out[1571][21]);
mul_8x8bit m4715 (image[621],filter[8],mul_out[1571][22]);

adder_8bit ad523 (mul_out[1569][20],mul_out[1569][21],mul_out[1569][22],mul_out[1570][20],mul_out[1570][21],mul_out[1570][22],mul_out[1571][20],mul_out[1571][21],mul_out[1571][22],conv_out[523]);



mul_8x8bit m4716 (image[564],filter[0],mul_out[1572][20]);
mul_8x8bit m4717 (image[565],filter[1],mul_out[1572][21]);
mul_8x8bit m4718 (image[566],filter[2],mul_out[1572][22]);
mul_8x8bit m4719 (image[592],filter[3],mul_out[1573][20]);
mul_8x8bit m4720 (image[593],filter[4],mul_out[1573][21]);
mul_8x8bit m4721 (image[594],filter[5],mul_out[1573][22]);
mul_8x8bit m4722 (image[620],filter[6],mul_out[1574][20]);
mul_8x8bit m4723 (image[621],filter[7],mul_out[1574][21]);
mul_8x8bit m4724 (image[622],filter[8],mul_out[1574][22]);

adder_8bit ad524 (mul_out[1572][20],mul_out[1572][21],mul_out[1572][22],mul_out[1573][20],mul_out[1573][21],mul_out[1573][22],mul_out[1574][20],mul_out[1574][21],mul_out[1574][22],conv_out[524]);



mul_8x8bit m4725 (image[565],filter[0],mul_out[1575][20]);
mul_8x8bit m4726 (image[566],filter[1],mul_out[1575][21]);
mul_8x8bit m4727 (image[567],filter[2],mul_out[1575][22]);
mul_8x8bit m4728 (image[593],filter[3],mul_out[1576][20]);
mul_8x8bit m4729 (image[594],filter[4],mul_out[1576][21]);
mul_8x8bit m4730 (image[595],filter[5],mul_out[1576][22]);
mul_8x8bit m4731 (image[621],filter[6],mul_out[1577][20]);
mul_8x8bit m4732 (image[622],filter[7],mul_out[1577][21]);
mul_8x8bit m4733 (image[623],filter[8],mul_out[1577][22]);

adder_8bit ad525 (mul_out[1575][20],mul_out[1575][21],mul_out[1575][22],mul_out[1576][20],mul_out[1576][21],mul_out[1576][22],mul_out[1577][20],mul_out[1577][21],mul_out[1577][22],conv_out[525]);



mul_8x8bit m4734 (image[566],filter[0],mul_out[1578][20]);
mul_8x8bit m4735 (image[567],filter[1],mul_out[1578][21]);
mul_8x8bit m4736 (image[568],filter[2],mul_out[1578][22]);
mul_8x8bit m4737 (image[594],filter[3],mul_out[1579][20]);
mul_8x8bit m4738 (image[595],filter[4],mul_out[1579][21]);
mul_8x8bit m4739 (image[596],filter[5],mul_out[1579][22]);
mul_8x8bit m4740 (image[622],filter[6],mul_out[1580][20]);
mul_8x8bit m4741 (image[623],filter[7],mul_out[1580][21]);
mul_8x8bit m4742 (image[624],filter[8],mul_out[1580][22]);

adder_8bit ad526 (mul_out[1578][20],mul_out[1578][21],mul_out[1578][22],mul_out[1579][20],mul_out[1579][21],mul_out[1579][22],mul_out[1580][20],mul_out[1580][21],mul_out[1580][22],conv_out[526]);



mul_8x8bit m4743 (image[567],filter[0],mul_out[1581][20]);
mul_8x8bit m4744 (image[568],filter[1],mul_out[1581][21]);
mul_8x8bit m4745 (image[569],filter[2],mul_out[1581][22]);
mul_8x8bit m4746 (image[595],filter[3],mul_out[1582][20]);
mul_8x8bit m4747 (image[596],filter[4],mul_out[1582][21]);
mul_8x8bit m4748 (image[597],filter[5],mul_out[1582][22]);
mul_8x8bit m4749 (image[623],filter[6],mul_out[1583][20]);
mul_8x8bit m4750 (image[624],filter[7],mul_out[1583][21]);
mul_8x8bit m4751 (image[625],filter[8],mul_out[1583][22]);

adder_8bit ad527 (mul_out[1581][20],mul_out[1581][21],mul_out[1581][22],mul_out[1582][20],mul_out[1582][21],mul_out[1582][22],mul_out[1583][20],mul_out[1583][21],mul_out[1583][22],conv_out[527]);



mul_8x8bit m4752 (image[568],filter[0],mul_out[1584][20]);
mul_8x8bit m4753 (image[569],filter[1],mul_out[1584][21]);
mul_8x8bit m4754 (image[570],filter[2],mul_out[1584][22]);
mul_8x8bit m4755 (image[596],filter[3],mul_out[1585][20]);
mul_8x8bit m4756 (image[597],filter[4],mul_out[1585][21]);
mul_8x8bit m4757 (image[598],filter[5],mul_out[1585][22]);
mul_8x8bit m4758 (image[624],filter[6],mul_out[1586][20]);
mul_8x8bit m4759 (image[625],filter[7],mul_out[1586][21]);
mul_8x8bit m4760 (image[626],filter[8],mul_out[1586][22]);

adder_8bit ad528 (mul_out[1584][20],mul_out[1584][21],mul_out[1584][22],mul_out[1585][20],mul_out[1585][21],mul_out[1585][22],mul_out[1586][20],mul_out[1586][21],mul_out[1586][22],conv_out[528]);



mul_8x8bit m4761 (image[569],filter[0],mul_out[1587][20]);
mul_8x8bit m4762 (image[570],filter[1],mul_out[1587][21]);
mul_8x8bit m4763 (image[571],filter[2],mul_out[1587][22]);
mul_8x8bit m4764 (image[597],filter[3],mul_out[1588][20]);
mul_8x8bit m4765 (image[598],filter[4],mul_out[1588][21]);
mul_8x8bit m4766 (image[599],filter[5],mul_out[1588][22]);
mul_8x8bit m4767 (image[625],filter[6],mul_out[1589][20]);
mul_8x8bit m4768 (image[626],filter[7],mul_out[1589][21]);
mul_8x8bit m4769 (image[627],filter[8],mul_out[1589][22]);

adder_8bit ad529 (mul_out[1587][20],mul_out[1587][21],mul_out[1587][22],mul_out[1588][20],mul_out[1588][21],mul_out[1588][22],mul_out[1589][20],mul_out[1589][21],mul_out[1589][22],conv_out[529]);



mul_8x8bit m4770 (image[570],filter[0],mul_out[1590][20]);
mul_8x8bit m4771 (image[571],filter[1],mul_out[1590][21]);
mul_8x8bit m4772 (image[572],filter[2],mul_out[1590][22]);
mul_8x8bit m4773 (image[598],filter[3],mul_out[1591][20]);
mul_8x8bit m4774 (image[599],filter[4],mul_out[1591][21]);
mul_8x8bit m4775 (image[600],filter[5],mul_out[1591][22]);
mul_8x8bit m4776 (image[626],filter[6],mul_out[1592][20]);
mul_8x8bit m4777 (image[627],filter[7],mul_out[1592][21]);
mul_8x8bit m4778 (image[628],filter[8],mul_out[1592][22]);

adder_8bit ad530 (mul_out[1590][20],mul_out[1590][21],mul_out[1590][22],mul_out[1591][20],mul_out[1591][21],mul_out[1591][22],mul_out[1592][20],mul_out[1592][21],mul_out[1592][22],conv_out[530]);



mul_8x8bit m4779 (image[571],filter[0],mul_out[1593][20]);
mul_8x8bit m4780 (image[572],filter[1],mul_out[1593][21]);
mul_8x8bit m4781 (image[573],filter[2],mul_out[1593][22]);
mul_8x8bit m4782 (image[599],filter[3],mul_out[1594][20]);
mul_8x8bit m4783 (image[600],filter[4],mul_out[1594][21]);
mul_8x8bit m4784 (image[601],filter[5],mul_out[1594][22]);
mul_8x8bit m4785 (image[627],filter[6],mul_out[1595][20]);
mul_8x8bit m4786 (image[628],filter[7],mul_out[1595][21]);
mul_8x8bit m4787 (image[629],filter[8],mul_out[1595][22]);

adder_8bit ad531 (mul_out[1593][20],mul_out[1593][21],mul_out[1593][22],mul_out[1594][20],mul_out[1594][21],mul_out[1594][22],mul_out[1595][20],mul_out[1595][21],mul_out[1595][22],conv_out[531]);



mul_8x8bit m4788 (image[572],filter[0],mul_out[1596][20]);
mul_8x8bit m4789 (image[573],filter[1],mul_out[1596][21]);
mul_8x8bit m4790 (image[574],filter[2],mul_out[1596][22]);
mul_8x8bit m4791 (image[600],filter[3],mul_out[1597][20]);
mul_8x8bit m4792 (image[601],filter[4],mul_out[1597][21]);
mul_8x8bit m4793 (image[602],filter[5],mul_out[1597][22]);
mul_8x8bit m4794 (image[628],filter[6],mul_out[1598][20]);
mul_8x8bit m4795 (image[629],filter[7],mul_out[1598][21]);
mul_8x8bit m4796 (image[630],filter[8],mul_out[1598][22]);

adder_8bit ad532 (mul_out[1596][20],mul_out[1596][21],mul_out[1596][22],mul_out[1597][20],mul_out[1597][21],mul_out[1597][22],mul_out[1598][20],mul_out[1598][21],mul_out[1598][22],conv_out[532]);



mul_8x8bit m4797 (image[573],filter[0],mul_out[1599][20]);
mul_8x8bit m4798 (image[574],filter[1],mul_out[1599][21]);
mul_8x8bit m4799 (image[575],filter[2],mul_out[1599][22]);
mul_8x8bit m4800 (image[601],filter[3],mul_out[1600][20]);
mul_8x8bit m4801 (image[602],filter[4],mul_out[1600][21]);
mul_8x8bit m4802 (image[603],filter[5],mul_out[1600][22]);
mul_8x8bit m4803 (image[629],filter[6],mul_out[1601][20]);
mul_8x8bit m4804 (image[630],filter[7],mul_out[1601][21]);
mul_8x8bit m4805 (image[631],filter[8],mul_out[1601][22]);

adder_8bit ad533 (mul_out[1599][20],mul_out[1599][21],mul_out[1599][22],mul_out[1600][20],mul_out[1600][21],mul_out[1600][22],mul_out[1601][20],mul_out[1601][21],mul_out[1601][22],conv_out[533]);



mul_8x8bit m4806 (image[574],filter[0],mul_out[1602][20]);
mul_8x8bit m4807 (image[575],filter[1],mul_out[1602][21]);
mul_8x8bit m4808 (image[576],filter[2],mul_out[1602][22]);
mul_8x8bit m4809 (image[602],filter[3],mul_out[1603][20]);
mul_8x8bit m4810 (image[603],filter[4],mul_out[1603][21]);
mul_8x8bit m4811 (image[604],filter[5],mul_out[1603][22]);
mul_8x8bit m4812 (image[630],filter[6],mul_out[1604][20]);
mul_8x8bit m4813 (image[631],filter[7],mul_out[1604][21]);
mul_8x8bit m4814 (image[632],filter[8],mul_out[1604][22]);

adder_8bit ad534 (mul_out[1602][20],mul_out[1602][21],mul_out[1602][22],mul_out[1603][20],mul_out[1603][21],mul_out[1603][22],mul_out[1604][20],mul_out[1604][21],mul_out[1604][22],conv_out[534]);



mul_8x8bit m4815 (image[575],filter[0],mul_out[1605][20]);
mul_8x8bit m4816 (image[576],filter[1],mul_out[1605][21]);
mul_8x8bit m4817 (image[577],filter[2],mul_out[1605][22]);
mul_8x8bit m4818 (image[603],filter[3],mul_out[1606][20]);
mul_8x8bit m4819 (image[604],filter[4],mul_out[1606][21]);
mul_8x8bit m4820 (image[605],filter[5],mul_out[1606][22]);
mul_8x8bit m4821 (image[631],filter[6],mul_out[1607][20]);
mul_8x8bit m4822 (image[632],filter[7],mul_out[1607][21]);
mul_8x8bit m4823 (image[633],filter[8],mul_out[1607][22]);

adder_8bit ad535 (mul_out[1605][20],mul_out[1605][21],mul_out[1605][22],mul_out[1606][20],mul_out[1606][21],mul_out[1606][22],mul_out[1607][20],mul_out[1607][21],mul_out[1607][22],conv_out[535]);



mul_8x8bit m4824 (image[576],filter[0],mul_out[1608][20]);
mul_8x8bit m4825 (image[577],filter[1],mul_out[1608][21]);
mul_8x8bit m4826 (image[578],filter[2],mul_out[1608][22]);
mul_8x8bit m4827 (image[604],filter[3],mul_out[1609][20]);
mul_8x8bit m4828 (image[605],filter[4],mul_out[1609][21]);
mul_8x8bit m4829 (image[606],filter[5],mul_out[1609][22]);
mul_8x8bit m4830 (image[632],filter[6],mul_out[1610][20]);
mul_8x8bit m4831 (image[633],filter[7],mul_out[1610][21]);
mul_8x8bit m4832 (image[634],filter[8],mul_out[1610][22]);

adder_8bit ad536 (mul_out[1608][20],mul_out[1608][21],mul_out[1608][22],mul_out[1609][20],mul_out[1609][21],mul_out[1609][22],mul_out[1610][20],mul_out[1610][21],mul_out[1610][22],conv_out[536]);



mul_8x8bit m4833 (image[577],filter[0],mul_out[1611][20]);
mul_8x8bit m4834 (image[578],filter[1],mul_out[1611][21]);
mul_8x8bit m4835 (image[579],filter[2],mul_out[1611][22]);
mul_8x8bit m4836 (image[605],filter[3],mul_out[1612][20]);
mul_8x8bit m4837 (image[606],filter[4],mul_out[1612][21]);
mul_8x8bit m4838 (image[607],filter[5],mul_out[1612][22]);
mul_8x8bit m4839 (image[633],filter[6],mul_out[1613][20]);
mul_8x8bit m4840 (image[634],filter[7],mul_out[1613][21]);
mul_8x8bit m4841 (image[635],filter[8],mul_out[1613][22]);

adder_8bit ad537 (mul_out[1611][20],mul_out[1611][21],mul_out[1611][22],mul_out[1612][20],mul_out[1612][21],mul_out[1612][22],mul_out[1613][20],mul_out[1613][21],mul_out[1613][22],conv_out[537]);



mul_8x8bit m4842 (image[578],filter[0],mul_out[1614][20]);
mul_8x8bit m4843 (image[579],filter[1],mul_out[1614][21]);
mul_8x8bit m4844 (image[580],filter[2],mul_out[1614][22]);
mul_8x8bit m4845 (image[606],filter[3],mul_out[1615][20]);
mul_8x8bit m4846 (image[607],filter[4],mul_out[1615][21]);
mul_8x8bit m4847 (image[608],filter[5],mul_out[1615][22]);
mul_8x8bit m4848 (image[634],filter[6],mul_out[1616][20]);
mul_8x8bit m4849 (image[635],filter[7],mul_out[1616][21]);
mul_8x8bit m4850 (image[636],filter[8],mul_out[1616][22]);

adder_8bit ad538 (mul_out[1614][20],mul_out[1614][21],mul_out[1614][22],mul_out[1615][20],mul_out[1615][21],mul_out[1615][22],mul_out[1616][20],mul_out[1616][21],mul_out[1616][22],conv_out[538]);



mul_8x8bit m4851 (image[579],filter[0],mul_out[1617][20]);
mul_8x8bit m4852 (image[580],filter[1],mul_out[1617][21]);
mul_8x8bit m4853 (image[581],filter[2],mul_out[1617][22]);
mul_8x8bit m4854 (image[607],filter[3],mul_out[1618][20]);
mul_8x8bit m4855 (image[608],filter[4],mul_out[1618][21]);
mul_8x8bit m4856 (image[609],filter[5],mul_out[1618][22]);
mul_8x8bit m4857 (image[635],filter[6],mul_out[1619][20]);
mul_8x8bit m4858 (image[636],filter[7],mul_out[1619][21]);
mul_8x8bit m4859 (image[637],filter[8],mul_out[1619][22]);

adder_8bit ad539 (mul_out[1617][20],mul_out[1617][21],mul_out[1617][22],mul_out[1618][20],mul_out[1618][21],mul_out[1618][22],mul_out[1619][20],mul_out[1619][21],mul_out[1619][22],conv_out[539]);



mul_8x8bit m4860 (image[580],filter[0],mul_out[1620][20]);
mul_8x8bit m4861 (image[581],filter[1],mul_out[1620][21]);
mul_8x8bit m4862 (image[582],filter[2],mul_out[1620][22]);
mul_8x8bit m4863 (image[608],filter[3],mul_out[1621][20]);
mul_8x8bit m4864 (image[609],filter[4],mul_out[1621][21]);
mul_8x8bit m4865 (image[610],filter[5],mul_out[1621][22]);
mul_8x8bit m4866 (image[636],filter[6],mul_out[1622][20]);
mul_8x8bit m4867 (image[637],filter[7],mul_out[1622][21]);
mul_8x8bit m4868 (image[638],filter[8],mul_out[1622][22]);

adder_8bit ad540 (mul_out[1620][20],mul_out[1620][21],mul_out[1620][22],mul_out[1621][20],mul_out[1621][21],mul_out[1621][22],mul_out[1622][20],mul_out[1622][21],mul_out[1622][22],conv_out[540]);



mul_8x8bit m4869 (image[581],filter[0],mul_out[1623][20]);
mul_8x8bit m4870 (image[582],filter[1],mul_out[1623][21]);
mul_8x8bit m4871 (image[583],filter[2],mul_out[1623][22]);
mul_8x8bit m4872 (image[609],filter[3],mul_out[1624][20]);
mul_8x8bit m4873 (image[610],filter[4],mul_out[1624][21]);
mul_8x8bit m4874 (image[611],filter[5],mul_out[1624][22]);
mul_8x8bit m4875 (image[637],filter[6],mul_out[1625][20]);
mul_8x8bit m4876 (image[638],filter[7],mul_out[1625][21]);
mul_8x8bit m4877 (image[639],filter[8],mul_out[1625][22]);

adder_8bit ad541 (mul_out[1623][20],mul_out[1623][21],mul_out[1623][22],mul_out[1624][20],mul_out[1624][21],mul_out[1624][22],mul_out[1625][20],mul_out[1625][21],mul_out[1625][22],conv_out[541]);



mul_8x8bit m4878 (image[582],filter[0],mul_out[1626][20]);
mul_8x8bit m4879 (image[583],filter[1],mul_out[1626][21]);
mul_8x8bit m4880 (image[584],filter[2],mul_out[1626][22]);
mul_8x8bit m4881 (image[610],filter[3],mul_out[1627][20]);
mul_8x8bit m4882 (image[611],filter[4],mul_out[1627][21]);
mul_8x8bit m4883 (image[612],filter[5],mul_out[1627][22]);
mul_8x8bit m4884 (image[638],filter[6],mul_out[1628][20]);
mul_8x8bit m4885 (image[639],filter[7],mul_out[1628][21]);
mul_8x8bit m4886 (image[640],filter[8],mul_out[1628][22]);

adder_8bit ad542 (mul_out[1626][20],mul_out[1626][21],mul_out[1626][22],mul_out[1627][20],mul_out[1627][21],mul_out[1627][22],mul_out[1628][20],mul_out[1628][21],mul_out[1628][22],conv_out[542]);



mul_8x8bit m4887 (image[583],filter[0],mul_out[1629][20]);
mul_8x8bit m4888 (image[584],filter[1],mul_out[1629][21]);
mul_8x8bit m4889 (image[585],filter[2],mul_out[1629][22]);
mul_8x8bit m4890 (image[611],filter[3],mul_out[1630][20]);
mul_8x8bit m4891 (image[612],filter[4],mul_out[1630][21]);
mul_8x8bit m4892 (image[613],filter[5],mul_out[1630][22]);
mul_8x8bit m4893 (image[639],filter[6],mul_out[1631][20]);
mul_8x8bit m4894 (image[640],filter[7],mul_out[1631][21]);
mul_8x8bit m4895 (image[641],filter[8],mul_out[1631][22]);

adder_8bit ad543 (mul_out[1629][20],mul_out[1629][21],mul_out[1629][22],mul_out[1630][20],mul_out[1630][21],mul_out[1630][22],mul_out[1631][20],mul_out[1631][21],mul_out[1631][22],conv_out[543]);



mul_8x8bit m4896 (image[584],filter[0],mul_out[1632][20]);
mul_8x8bit m4897 (image[585],filter[1],mul_out[1632][21]);
mul_8x8bit m4898 (image[586],filter[2],mul_out[1632][22]);
mul_8x8bit m4899 (image[612],filter[3],mul_out[1633][20]);
mul_8x8bit m4900 (image[613],filter[4],mul_out[1633][21]);
mul_8x8bit m4901 (image[614],filter[5],mul_out[1633][22]);
mul_8x8bit m4902 (image[640],filter[6],mul_out[1634][20]);
mul_8x8bit m4903 (image[641],filter[7],mul_out[1634][21]);
mul_8x8bit m4904 (image[642],filter[8],mul_out[1634][22]);

adder_8bit ad544 (mul_out[1632][20],mul_out[1632][21],mul_out[1632][22],mul_out[1633][20],mul_out[1633][21],mul_out[1633][22],mul_out[1634][20],mul_out[1634][21],mul_out[1634][22],conv_out[544]);



mul_8x8bit m4905 (image[585],filter[0],mul_out[1635][20]);
mul_8x8bit m4906 (image[586],filter[1],mul_out[1635][21]);
mul_8x8bit m4907 (image[587],filter[2],mul_out[1635][22]);
mul_8x8bit m4908 (image[613],filter[3],mul_out[1636][20]);
mul_8x8bit m4909 (image[614],filter[4],mul_out[1636][21]);
mul_8x8bit m4910 (image[615],filter[5],mul_out[1636][22]);
mul_8x8bit m4911 (image[641],filter[6],mul_out[1637][20]);
mul_8x8bit m4912 (image[642],filter[7],mul_out[1637][21]);
mul_8x8bit m4913 (image[643],filter[8],mul_out[1637][22]);

adder_8bit ad545 (mul_out[1635][20],mul_out[1635][21],mul_out[1635][22],mul_out[1636][20],mul_out[1636][21],mul_out[1636][22],mul_out[1637][20],mul_out[1637][21],mul_out[1637][22],conv_out[545]);



mul_8x8bit m4914 (image[588],filter[0],mul_out[1638][21]);
mul_8x8bit m4915 (image[589],filter[1],mul_out[1638][22]);
mul_8x8bit m4916 (image[590],filter[2],mul_out[1638][23]);
mul_8x8bit m4917 (image[616],filter[3],mul_out[1639][21]);
mul_8x8bit m4918 (image[617],filter[4],mul_out[1639][22]);
mul_8x8bit m4919 (image[618],filter[5],mul_out[1639][23]);
mul_8x8bit m4920 (image[644],filter[6],mul_out[1640][21]);
mul_8x8bit m4921 (image[645],filter[7],mul_out[1640][22]);
mul_8x8bit m4922 (image[646],filter[8],mul_out[1640][23]);

adder_8bit ad546 (mul_out[1638][21],mul_out[1638][22],mul_out[1638][23],mul_out[1639][21],mul_out[1639][22],mul_out[1639][23],mul_out[1640][21],mul_out[1640][22],mul_out[1640][23],conv_out[546]);



mul_8x8bit m4923 (image[589],filter[0],mul_out[1641][21]);
mul_8x8bit m4924 (image[590],filter[1],mul_out[1641][22]);
mul_8x8bit m4925 (image[591],filter[2],mul_out[1641][23]);
mul_8x8bit m4926 (image[617],filter[3],mul_out[1642][21]);
mul_8x8bit m4927 (image[618],filter[4],mul_out[1642][22]);
mul_8x8bit m4928 (image[619],filter[5],mul_out[1642][23]);
mul_8x8bit m4929 (image[645],filter[6],mul_out[1643][21]);
mul_8x8bit m4930 (image[646],filter[7],mul_out[1643][22]);
mul_8x8bit m4931 (image[647],filter[8],mul_out[1643][23]);

adder_8bit ad547 (mul_out[1641][21],mul_out[1641][22],mul_out[1641][23],mul_out[1642][21],mul_out[1642][22],mul_out[1642][23],mul_out[1643][21],mul_out[1643][22],mul_out[1643][23],conv_out[547]);



mul_8x8bit m4932 (image[590],filter[0],mul_out[1644][21]);
mul_8x8bit m4933 (image[591],filter[1],mul_out[1644][22]);
mul_8x8bit m4934 (image[592],filter[2],mul_out[1644][23]);
mul_8x8bit m4935 (image[618],filter[3],mul_out[1645][21]);
mul_8x8bit m4936 (image[619],filter[4],mul_out[1645][22]);
mul_8x8bit m4937 (image[620],filter[5],mul_out[1645][23]);
mul_8x8bit m4938 (image[646],filter[6],mul_out[1646][21]);
mul_8x8bit m4939 (image[647],filter[7],mul_out[1646][22]);
mul_8x8bit m4940 (image[648],filter[8],mul_out[1646][23]);

adder_8bit ad548 (mul_out[1644][21],mul_out[1644][22],mul_out[1644][23],mul_out[1645][21],mul_out[1645][22],mul_out[1645][23],mul_out[1646][21],mul_out[1646][22],mul_out[1646][23],conv_out[548]);



mul_8x8bit m4941 (image[591],filter[0],mul_out[1647][21]);
mul_8x8bit m4942 (image[592],filter[1],mul_out[1647][22]);
mul_8x8bit m4943 (image[593],filter[2],mul_out[1647][23]);
mul_8x8bit m4944 (image[619],filter[3],mul_out[1648][21]);
mul_8x8bit m4945 (image[620],filter[4],mul_out[1648][22]);
mul_8x8bit m4946 (image[621],filter[5],mul_out[1648][23]);
mul_8x8bit m4947 (image[647],filter[6],mul_out[1649][21]);
mul_8x8bit m4948 (image[648],filter[7],mul_out[1649][22]);
mul_8x8bit m4949 (image[649],filter[8],mul_out[1649][23]);

adder_8bit ad549 (mul_out[1647][21],mul_out[1647][22],mul_out[1647][23],mul_out[1648][21],mul_out[1648][22],mul_out[1648][23],mul_out[1649][21],mul_out[1649][22],mul_out[1649][23],conv_out[549]);



mul_8x8bit m4950 (image[592],filter[0],mul_out[1650][21]);
mul_8x8bit m4951 (image[593],filter[1],mul_out[1650][22]);
mul_8x8bit m4952 (image[594],filter[2],mul_out[1650][23]);
mul_8x8bit m4953 (image[620],filter[3],mul_out[1651][21]);
mul_8x8bit m4954 (image[621],filter[4],mul_out[1651][22]);
mul_8x8bit m4955 (image[622],filter[5],mul_out[1651][23]);
mul_8x8bit m4956 (image[648],filter[6],mul_out[1652][21]);
mul_8x8bit m4957 (image[649],filter[7],mul_out[1652][22]);
mul_8x8bit m4958 (image[650],filter[8],mul_out[1652][23]);

adder_8bit ad550 (mul_out[1650][21],mul_out[1650][22],mul_out[1650][23],mul_out[1651][21],mul_out[1651][22],mul_out[1651][23],mul_out[1652][21],mul_out[1652][22],mul_out[1652][23],conv_out[550]);



mul_8x8bit m4959 (image[593],filter[0],mul_out[1653][21]);
mul_8x8bit m4960 (image[594],filter[1],mul_out[1653][22]);
mul_8x8bit m4961 (image[595],filter[2],mul_out[1653][23]);
mul_8x8bit m4962 (image[621],filter[3],mul_out[1654][21]);
mul_8x8bit m4963 (image[622],filter[4],mul_out[1654][22]);
mul_8x8bit m4964 (image[623],filter[5],mul_out[1654][23]);
mul_8x8bit m4965 (image[649],filter[6],mul_out[1655][21]);
mul_8x8bit m4966 (image[650],filter[7],mul_out[1655][22]);
mul_8x8bit m4967 (image[651],filter[8],mul_out[1655][23]);

adder_8bit ad551 (mul_out[1653][21],mul_out[1653][22],mul_out[1653][23],mul_out[1654][21],mul_out[1654][22],mul_out[1654][23],mul_out[1655][21],mul_out[1655][22],mul_out[1655][23],conv_out[551]);



mul_8x8bit m4968 (image[594],filter[0],mul_out[1656][21]);
mul_8x8bit m4969 (image[595],filter[1],mul_out[1656][22]);
mul_8x8bit m4970 (image[596],filter[2],mul_out[1656][23]);
mul_8x8bit m4971 (image[622],filter[3],mul_out[1657][21]);
mul_8x8bit m4972 (image[623],filter[4],mul_out[1657][22]);
mul_8x8bit m4973 (image[624],filter[5],mul_out[1657][23]);
mul_8x8bit m4974 (image[650],filter[6],mul_out[1658][21]);
mul_8x8bit m4975 (image[651],filter[7],mul_out[1658][22]);
mul_8x8bit m4976 (image[652],filter[8],mul_out[1658][23]);

adder_8bit ad552 (mul_out[1656][21],mul_out[1656][22],mul_out[1656][23],mul_out[1657][21],mul_out[1657][22],mul_out[1657][23],mul_out[1658][21],mul_out[1658][22],mul_out[1658][23],conv_out[552]);



mul_8x8bit m4977 (image[595],filter[0],mul_out[1659][21]);
mul_8x8bit m4978 (image[596],filter[1],mul_out[1659][22]);
mul_8x8bit m4979 (image[597],filter[2],mul_out[1659][23]);
mul_8x8bit m4980 (image[623],filter[3],mul_out[1660][21]);
mul_8x8bit m4981 (image[624],filter[4],mul_out[1660][22]);
mul_8x8bit m4982 (image[625],filter[5],mul_out[1660][23]);
mul_8x8bit m4983 (image[651],filter[6],mul_out[1661][21]);
mul_8x8bit m4984 (image[652],filter[7],mul_out[1661][22]);
mul_8x8bit m4985 (image[653],filter[8],mul_out[1661][23]);

adder_8bit ad553 (mul_out[1659][21],mul_out[1659][22],mul_out[1659][23],mul_out[1660][21],mul_out[1660][22],mul_out[1660][23],mul_out[1661][21],mul_out[1661][22],mul_out[1661][23],conv_out[553]);



mul_8x8bit m4986 (image[596],filter[0],mul_out[1662][21]);
mul_8x8bit m4987 (image[597],filter[1],mul_out[1662][22]);
mul_8x8bit m4988 (image[598],filter[2],mul_out[1662][23]);
mul_8x8bit m4989 (image[624],filter[3],mul_out[1663][21]);
mul_8x8bit m4990 (image[625],filter[4],mul_out[1663][22]);
mul_8x8bit m4991 (image[626],filter[5],mul_out[1663][23]);
mul_8x8bit m4992 (image[652],filter[6],mul_out[1664][21]);
mul_8x8bit m4993 (image[653],filter[7],mul_out[1664][22]);
mul_8x8bit m4994 (image[654],filter[8],mul_out[1664][23]);

adder_8bit ad554 (mul_out[1662][21],mul_out[1662][22],mul_out[1662][23],mul_out[1663][21],mul_out[1663][22],mul_out[1663][23],mul_out[1664][21],mul_out[1664][22],mul_out[1664][23],conv_out[554]);



mul_8x8bit m4995 (image[597],filter[0],mul_out[1665][21]);
mul_8x8bit m4996 (image[598],filter[1],mul_out[1665][22]);
mul_8x8bit m4997 (image[599],filter[2],mul_out[1665][23]);
mul_8x8bit m4998 (image[625],filter[3],mul_out[1666][21]);
mul_8x8bit m4999 (image[626],filter[4],mul_out[1666][22]);
mul_8x8bit m5000 (image[627],filter[5],mul_out[1666][23]);
mul_8x8bit m5001 (image[653],filter[6],mul_out[1667][21]);
mul_8x8bit m5002 (image[654],filter[7],mul_out[1667][22]);
mul_8x8bit m5003 (image[655],filter[8],mul_out[1667][23]);

adder_8bit ad555 (mul_out[1665][21],mul_out[1665][22],mul_out[1665][23],mul_out[1666][21],mul_out[1666][22],mul_out[1666][23],mul_out[1667][21],mul_out[1667][22],mul_out[1667][23],conv_out[555]);



mul_8x8bit m5004 (image[598],filter[0],mul_out[1668][21]);
mul_8x8bit m5005 (image[599],filter[1],mul_out[1668][22]);
mul_8x8bit m5006 (image[600],filter[2],mul_out[1668][23]);
mul_8x8bit m5007 (image[626],filter[3],mul_out[1669][21]);
mul_8x8bit m5008 (image[627],filter[4],mul_out[1669][22]);
mul_8x8bit m5009 (image[628],filter[5],mul_out[1669][23]);
mul_8x8bit m5010 (image[654],filter[6],mul_out[1670][21]);
mul_8x8bit m5011 (image[655],filter[7],mul_out[1670][22]);
mul_8x8bit m5012 (image[656],filter[8],mul_out[1670][23]);

adder_8bit ad556 (mul_out[1668][21],mul_out[1668][22],mul_out[1668][23],mul_out[1669][21],mul_out[1669][22],mul_out[1669][23],mul_out[1670][21],mul_out[1670][22],mul_out[1670][23],conv_out[556]);



mul_8x8bit m5013 (image[599],filter[0],mul_out[1671][21]);
mul_8x8bit m5014 (image[600],filter[1],mul_out[1671][22]);
mul_8x8bit m5015 (image[601],filter[2],mul_out[1671][23]);
mul_8x8bit m5016 (image[627],filter[3],mul_out[1672][21]);
mul_8x8bit m5017 (image[628],filter[4],mul_out[1672][22]);
mul_8x8bit m5018 (image[629],filter[5],mul_out[1672][23]);
mul_8x8bit m5019 (image[655],filter[6],mul_out[1673][21]);
mul_8x8bit m5020 (image[656],filter[7],mul_out[1673][22]);
mul_8x8bit m5021 (image[657],filter[8],mul_out[1673][23]);

adder_8bit ad557 (mul_out[1671][21],mul_out[1671][22],mul_out[1671][23],mul_out[1672][21],mul_out[1672][22],mul_out[1672][23],mul_out[1673][21],mul_out[1673][22],mul_out[1673][23],conv_out[557]);



mul_8x8bit m5022 (image[600],filter[0],mul_out[1674][21]);
mul_8x8bit m5023 (image[601],filter[1],mul_out[1674][22]);
mul_8x8bit m5024 (image[602],filter[2],mul_out[1674][23]);
mul_8x8bit m5025 (image[628],filter[3],mul_out[1675][21]);
mul_8x8bit m5026 (image[629],filter[4],mul_out[1675][22]);
mul_8x8bit m5027 (image[630],filter[5],mul_out[1675][23]);
mul_8x8bit m5028 (image[656],filter[6],mul_out[1676][21]);
mul_8x8bit m5029 (image[657],filter[7],mul_out[1676][22]);
mul_8x8bit m5030 (image[658],filter[8],mul_out[1676][23]);

adder_8bit ad558 (mul_out[1674][21],mul_out[1674][22],mul_out[1674][23],mul_out[1675][21],mul_out[1675][22],mul_out[1675][23],mul_out[1676][21],mul_out[1676][22],mul_out[1676][23],conv_out[558]);



mul_8x8bit m5031 (image[601],filter[0],mul_out[1677][21]);
mul_8x8bit m5032 (image[602],filter[1],mul_out[1677][22]);
mul_8x8bit m5033 (image[603],filter[2],mul_out[1677][23]);
mul_8x8bit m5034 (image[629],filter[3],mul_out[1678][21]);
mul_8x8bit m5035 (image[630],filter[4],mul_out[1678][22]);
mul_8x8bit m5036 (image[631],filter[5],mul_out[1678][23]);
mul_8x8bit m5037 (image[657],filter[6],mul_out[1679][21]);
mul_8x8bit m5038 (image[658],filter[7],mul_out[1679][22]);
mul_8x8bit m5039 (image[659],filter[8],mul_out[1679][23]);

adder_8bit ad559 (mul_out[1677][21],mul_out[1677][22],mul_out[1677][23],mul_out[1678][21],mul_out[1678][22],mul_out[1678][23],mul_out[1679][21],mul_out[1679][22],mul_out[1679][23],conv_out[559]);



mul_8x8bit m5040 (image[602],filter[0],mul_out[1680][21]);
mul_8x8bit m5041 (image[603],filter[1],mul_out[1680][22]);
mul_8x8bit m5042 (image[604],filter[2],mul_out[1680][23]);
mul_8x8bit m5043 (image[630],filter[3],mul_out[1681][21]);
mul_8x8bit m5044 (image[631],filter[4],mul_out[1681][22]);
mul_8x8bit m5045 (image[632],filter[5],mul_out[1681][23]);
mul_8x8bit m5046 (image[658],filter[6],mul_out[1682][21]);
mul_8x8bit m5047 (image[659],filter[7],mul_out[1682][22]);
mul_8x8bit m5048 (image[660],filter[8],mul_out[1682][23]);

adder_8bit ad560 (mul_out[1680][21],mul_out[1680][22],mul_out[1680][23],mul_out[1681][21],mul_out[1681][22],mul_out[1681][23],mul_out[1682][21],mul_out[1682][22],mul_out[1682][23],conv_out[560]);



mul_8x8bit m5049 (image[603],filter[0],mul_out[1683][21]);
mul_8x8bit m5050 (image[604],filter[1],mul_out[1683][22]);
mul_8x8bit m5051 (image[605],filter[2],mul_out[1683][23]);
mul_8x8bit m5052 (image[631],filter[3],mul_out[1684][21]);
mul_8x8bit m5053 (image[632],filter[4],mul_out[1684][22]);
mul_8x8bit m5054 (image[633],filter[5],mul_out[1684][23]);
mul_8x8bit m5055 (image[659],filter[6],mul_out[1685][21]);
mul_8x8bit m5056 (image[660],filter[7],mul_out[1685][22]);
mul_8x8bit m5057 (image[661],filter[8],mul_out[1685][23]);

adder_8bit ad561 (mul_out[1683][21],mul_out[1683][22],mul_out[1683][23],mul_out[1684][21],mul_out[1684][22],mul_out[1684][23],mul_out[1685][21],mul_out[1685][22],mul_out[1685][23],conv_out[561]);



mul_8x8bit m5058 (image[604],filter[0],mul_out[1686][21]);
mul_8x8bit m5059 (image[605],filter[1],mul_out[1686][22]);
mul_8x8bit m5060 (image[606],filter[2],mul_out[1686][23]);
mul_8x8bit m5061 (image[632],filter[3],mul_out[1687][21]);
mul_8x8bit m5062 (image[633],filter[4],mul_out[1687][22]);
mul_8x8bit m5063 (image[634],filter[5],mul_out[1687][23]);
mul_8x8bit m5064 (image[660],filter[6],mul_out[1688][21]);
mul_8x8bit m5065 (image[661],filter[7],mul_out[1688][22]);
mul_8x8bit m5066 (image[662],filter[8],mul_out[1688][23]);

adder_8bit ad562 (mul_out[1686][21],mul_out[1686][22],mul_out[1686][23],mul_out[1687][21],mul_out[1687][22],mul_out[1687][23],mul_out[1688][21],mul_out[1688][22],mul_out[1688][23],conv_out[562]);



mul_8x8bit m5067 (image[605],filter[0],mul_out[1689][21]);
mul_8x8bit m5068 (image[606],filter[1],mul_out[1689][22]);
mul_8x8bit m5069 (image[607],filter[2],mul_out[1689][23]);
mul_8x8bit m5070 (image[633],filter[3],mul_out[1690][21]);
mul_8x8bit m5071 (image[634],filter[4],mul_out[1690][22]);
mul_8x8bit m5072 (image[635],filter[5],mul_out[1690][23]);
mul_8x8bit m5073 (image[661],filter[6],mul_out[1691][21]);
mul_8x8bit m5074 (image[662],filter[7],mul_out[1691][22]);
mul_8x8bit m5075 (image[663],filter[8],mul_out[1691][23]);

adder_8bit ad563 (mul_out[1689][21],mul_out[1689][22],mul_out[1689][23],mul_out[1690][21],mul_out[1690][22],mul_out[1690][23],mul_out[1691][21],mul_out[1691][22],mul_out[1691][23],conv_out[563]);



mul_8x8bit m5076 (image[606],filter[0],mul_out[1692][21]);
mul_8x8bit m5077 (image[607],filter[1],mul_out[1692][22]);
mul_8x8bit m5078 (image[608],filter[2],mul_out[1692][23]);
mul_8x8bit m5079 (image[634],filter[3],mul_out[1693][21]);
mul_8x8bit m5080 (image[635],filter[4],mul_out[1693][22]);
mul_8x8bit m5081 (image[636],filter[5],mul_out[1693][23]);
mul_8x8bit m5082 (image[662],filter[6],mul_out[1694][21]);
mul_8x8bit m5083 (image[663],filter[7],mul_out[1694][22]);
mul_8x8bit m5084 (image[664],filter[8],mul_out[1694][23]);

adder_8bit ad564 (mul_out[1692][21],mul_out[1692][22],mul_out[1692][23],mul_out[1693][21],mul_out[1693][22],mul_out[1693][23],mul_out[1694][21],mul_out[1694][22],mul_out[1694][23],conv_out[564]);



mul_8x8bit m5085 (image[607],filter[0],mul_out[1695][21]);
mul_8x8bit m5086 (image[608],filter[1],mul_out[1695][22]);
mul_8x8bit m5087 (image[609],filter[2],mul_out[1695][23]);
mul_8x8bit m5088 (image[635],filter[3],mul_out[1696][21]);
mul_8x8bit m5089 (image[636],filter[4],mul_out[1696][22]);
mul_8x8bit m5090 (image[637],filter[5],mul_out[1696][23]);
mul_8x8bit m5091 (image[663],filter[6],mul_out[1697][21]);
mul_8x8bit m5092 (image[664],filter[7],mul_out[1697][22]);
mul_8x8bit m5093 (image[665],filter[8],mul_out[1697][23]);

adder_8bit ad565 (mul_out[1695][21],mul_out[1695][22],mul_out[1695][23],mul_out[1696][21],mul_out[1696][22],mul_out[1696][23],mul_out[1697][21],mul_out[1697][22],mul_out[1697][23],conv_out[565]);



mul_8x8bit m5094 (image[608],filter[0],mul_out[1698][21]);
mul_8x8bit m5095 (image[609],filter[1],mul_out[1698][22]);
mul_8x8bit m5096 (image[610],filter[2],mul_out[1698][23]);
mul_8x8bit m5097 (image[636],filter[3],mul_out[1699][21]);
mul_8x8bit m5098 (image[637],filter[4],mul_out[1699][22]);
mul_8x8bit m5099 (image[638],filter[5],mul_out[1699][23]);
mul_8x8bit m5100 (image[664],filter[6],mul_out[1700][21]);
mul_8x8bit m5101 (image[665],filter[7],mul_out[1700][22]);
mul_8x8bit m5102 (image[666],filter[8],mul_out[1700][23]);

adder_8bit ad566 (mul_out[1698][21],mul_out[1698][22],mul_out[1698][23],mul_out[1699][21],mul_out[1699][22],mul_out[1699][23],mul_out[1700][21],mul_out[1700][22],mul_out[1700][23],conv_out[566]);



mul_8x8bit m5103 (image[609],filter[0],mul_out[1701][21]);
mul_8x8bit m5104 (image[610],filter[1],mul_out[1701][22]);
mul_8x8bit m5105 (image[611],filter[2],mul_out[1701][23]);
mul_8x8bit m5106 (image[637],filter[3],mul_out[1702][21]);
mul_8x8bit m5107 (image[638],filter[4],mul_out[1702][22]);
mul_8x8bit m5108 (image[639],filter[5],mul_out[1702][23]);
mul_8x8bit m5109 (image[665],filter[6],mul_out[1703][21]);
mul_8x8bit m5110 (image[666],filter[7],mul_out[1703][22]);
mul_8x8bit m5111 (image[667],filter[8],mul_out[1703][23]);

adder_8bit ad567 (mul_out[1701][21],mul_out[1701][22],mul_out[1701][23],mul_out[1702][21],mul_out[1702][22],mul_out[1702][23],mul_out[1703][21],mul_out[1703][22],mul_out[1703][23],conv_out[567]);



mul_8x8bit m5112 (image[610],filter[0],mul_out[1704][21]);
mul_8x8bit m5113 (image[611],filter[1],mul_out[1704][22]);
mul_8x8bit m5114 (image[612],filter[2],mul_out[1704][23]);
mul_8x8bit m5115 (image[638],filter[3],mul_out[1705][21]);
mul_8x8bit m5116 (image[639],filter[4],mul_out[1705][22]);
mul_8x8bit m5117 (image[640],filter[5],mul_out[1705][23]);
mul_8x8bit m5118 (image[666],filter[6],mul_out[1706][21]);
mul_8x8bit m5119 (image[667],filter[7],mul_out[1706][22]);
mul_8x8bit m5120 (image[668],filter[8],mul_out[1706][23]);

adder_8bit ad568 (mul_out[1704][21],mul_out[1704][22],mul_out[1704][23],mul_out[1705][21],mul_out[1705][22],mul_out[1705][23],mul_out[1706][21],mul_out[1706][22],mul_out[1706][23],conv_out[568]);



mul_8x8bit m5121 (image[611],filter[0],mul_out[1707][21]);
mul_8x8bit m5122 (image[612],filter[1],mul_out[1707][22]);
mul_8x8bit m5123 (image[613],filter[2],mul_out[1707][23]);
mul_8x8bit m5124 (image[639],filter[3],mul_out[1708][21]);
mul_8x8bit m5125 (image[640],filter[4],mul_out[1708][22]);
mul_8x8bit m5126 (image[641],filter[5],mul_out[1708][23]);
mul_8x8bit m5127 (image[667],filter[6],mul_out[1709][21]);
mul_8x8bit m5128 (image[668],filter[7],mul_out[1709][22]);
mul_8x8bit m5129 (image[669],filter[8],mul_out[1709][23]);

adder_8bit ad569 (mul_out[1707][21],mul_out[1707][22],mul_out[1707][23],mul_out[1708][21],mul_out[1708][22],mul_out[1708][23],mul_out[1709][21],mul_out[1709][22],mul_out[1709][23],conv_out[569]);



mul_8x8bit m5130 (image[612],filter[0],mul_out[1710][21]);
mul_8x8bit m5131 (image[613],filter[1],mul_out[1710][22]);
mul_8x8bit m5132 (image[614],filter[2],mul_out[1710][23]);
mul_8x8bit m5133 (image[640],filter[3],mul_out[1711][21]);
mul_8x8bit m5134 (image[641],filter[4],mul_out[1711][22]);
mul_8x8bit m5135 (image[642],filter[5],mul_out[1711][23]);
mul_8x8bit m5136 (image[668],filter[6],mul_out[1712][21]);
mul_8x8bit m5137 (image[669],filter[7],mul_out[1712][22]);
mul_8x8bit m5138 (image[670],filter[8],mul_out[1712][23]);

adder_8bit ad570 (mul_out[1710][21],mul_out[1710][22],mul_out[1710][23],mul_out[1711][21],mul_out[1711][22],mul_out[1711][23],mul_out[1712][21],mul_out[1712][22],mul_out[1712][23],conv_out[570]);



mul_8x8bit m5139 (image[613],filter[0],mul_out[1713][21]);
mul_8x8bit m5140 (image[614],filter[1],mul_out[1713][22]);
mul_8x8bit m5141 (image[615],filter[2],mul_out[1713][23]);
mul_8x8bit m5142 (image[641],filter[3],mul_out[1714][21]);
mul_8x8bit m5143 (image[642],filter[4],mul_out[1714][22]);
mul_8x8bit m5144 (image[643],filter[5],mul_out[1714][23]);
mul_8x8bit m5145 (image[669],filter[6],mul_out[1715][21]);
mul_8x8bit m5146 (image[670],filter[7],mul_out[1715][22]);
mul_8x8bit m5147 (image[671],filter[8],mul_out[1715][23]);

adder_8bit ad571 (mul_out[1713][21],mul_out[1713][22],mul_out[1713][23],mul_out[1714][21],mul_out[1714][22],mul_out[1714][23],mul_out[1715][21],mul_out[1715][22],mul_out[1715][23],conv_out[571]);



mul_8x8bit m5148 (image[616],filter[0],mul_out[1716][22]);
mul_8x8bit m5149 (image[617],filter[1],mul_out[1716][23]);
mul_8x8bit m5150 (image[618],filter[2],mul_out[1716][24]);
mul_8x8bit m5151 (image[644],filter[3],mul_out[1717][22]);
mul_8x8bit m5152 (image[645],filter[4],mul_out[1717][23]);
mul_8x8bit m5153 (image[646],filter[5],mul_out[1717][24]);
mul_8x8bit m5154 (image[672],filter[6],mul_out[1718][22]);
mul_8x8bit m5155 (image[673],filter[7],mul_out[1718][23]);
mul_8x8bit m5156 (image[674],filter[8],mul_out[1718][24]);

adder_8bit ad572 (mul_out[1716][22],mul_out[1716][23],mul_out[1716][24],mul_out[1717][22],mul_out[1717][23],mul_out[1717][24],mul_out[1718][22],mul_out[1718][23],mul_out[1718][24],conv_out[572]);



mul_8x8bit m5157 (image[617],filter[0],mul_out[1719][22]);
mul_8x8bit m5158 (image[618],filter[1],mul_out[1719][23]);
mul_8x8bit m5159 (image[619],filter[2],mul_out[1719][24]);
mul_8x8bit m5160 (image[645],filter[3],mul_out[1720][22]);
mul_8x8bit m5161 (image[646],filter[4],mul_out[1720][23]);
mul_8x8bit m5162 (image[647],filter[5],mul_out[1720][24]);
mul_8x8bit m5163 (image[673],filter[6],mul_out[1721][22]);
mul_8x8bit m5164 (image[674],filter[7],mul_out[1721][23]);
mul_8x8bit m5165 (image[675],filter[8],mul_out[1721][24]);

adder_8bit ad573 (mul_out[1719][22],mul_out[1719][23],mul_out[1719][24],mul_out[1720][22],mul_out[1720][23],mul_out[1720][24],mul_out[1721][22],mul_out[1721][23],mul_out[1721][24],conv_out[573]);



mul_8x8bit m5166 (image[618],filter[0],mul_out[1722][22]);
mul_8x8bit m5167 (image[619],filter[1],mul_out[1722][23]);
mul_8x8bit m5168 (image[620],filter[2],mul_out[1722][24]);
mul_8x8bit m5169 (image[646],filter[3],mul_out[1723][22]);
mul_8x8bit m5170 (image[647],filter[4],mul_out[1723][23]);
mul_8x8bit m5171 (image[648],filter[5],mul_out[1723][24]);
mul_8x8bit m5172 (image[674],filter[6],mul_out[1724][22]);
mul_8x8bit m5173 (image[675],filter[7],mul_out[1724][23]);
mul_8x8bit m5174 (image[676],filter[8],mul_out[1724][24]);

adder_8bit ad574 (mul_out[1722][22],mul_out[1722][23],mul_out[1722][24],mul_out[1723][22],mul_out[1723][23],mul_out[1723][24],mul_out[1724][22],mul_out[1724][23],mul_out[1724][24],conv_out[574]);



mul_8x8bit m5175 (image[619],filter[0],mul_out[1725][22]);
mul_8x8bit m5176 (image[620],filter[1],mul_out[1725][23]);
mul_8x8bit m5177 (image[621],filter[2],mul_out[1725][24]);
mul_8x8bit m5178 (image[647],filter[3],mul_out[1726][22]);
mul_8x8bit m5179 (image[648],filter[4],mul_out[1726][23]);
mul_8x8bit m5180 (image[649],filter[5],mul_out[1726][24]);
mul_8x8bit m5181 (image[675],filter[6],mul_out[1727][22]);
mul_8x8bit m5182 (image[676],filter[7],mul_out[1727][23]);
mul_8x8bit m5183 (image[677],filter[8],mul_out[1727][24]);

adder_8bit ad575 (mul_out[1725][22],mul_out[1725][23],mul_out[1725][24],mul_out[1726][22],mul_out[1726][23],mul_out[1726][24],mul_out[1727][22],mul_out[1727][23],mul_out[1727][24],conv_out[575]);



mul_8x8bit m5184 (image[620],filter[0],mul_out[1728][22]);
mul_8x8bit m5185 (image[621],filter[1],mul_out[1728][23]);
mul_8x8bit m5186 (image[622],filter[2],mul_out[1728][24]);
mul_8x8bit m5187 (image[648],filter[3],mul_out[1729][22]);
mul_8x8bit m5188 (image[649],filter[4],mul_out[1729][23]);
mul_8x8bit m5189 (image[650],filter[5],mul_out[1729][24]);
mul_8x8bit m5190 (image[676],filter[6],mul_out[1730][22]);
mul_8x8bit m5191 (image[677],filter[7],mul_out[1730][23]);
mul_8x8bit m5192 (image[678],filter[8],mul_out[1730][24]);

adder_8bit ad576 (mul_out[1728][22],mul_out[1728][23],mul_out[1728][24],mul_out[1729][22],mul_out[1729][23],mul_out[1729][24],mul_out[1730][22],mul_out[1730][23],mul_out[1730][24],conv_out[576]);



mul_8x8bit m5193 (image[621],filter[0],mul_out[1731][22]);
mul_8x8bit m5194 (image[622],filter[1],mul_out[1731][23]);
mul_8x8bit m5195 (image[623],filter[2],mul_out[1731][24]);
mul_8x8bit m5196 (image[649],filter[3],mul_out[1732][22]);
mul_8x8bit m5197 (image[650],filter[4],mul_out[1732][23]);
mul_8x8bit m5198 (image[651],filter[5],mul_out[1732][24]);
mul_8x8bit m5199 (image[677],filter[6],mul_out[1733][22]);
mul_8x8bit m5200 (image[678],filter[7],mul_out[1733][23]);
mul_8x8bit m5201 (image[679],filter[8],mul_out[1733][24]);

adder_8bit ad577 (mul_out[1731][22],mul_out[1731][23],mul_out[1731][24],mul_out[1732][22],mul_out[1732][23],mul_out[1732][24],mul_out[1733][22],mul_out[1733][23],mul_out[1733][24],conv_out[577]);



mul_8x8bit m5202 (image[622],filter[0],mul_out[1734][22]);
mul_8x8bit m5203 (image[623],filter[1],mul_out[1734][23]);
mul_8x8bit m5204 (image[624],filter[2],mul_out[1734][24]);
mul_8x8bit m5205 (image[650],filter[3],mul_out[1735][22]);
mul_8x8bit m5206 (image[651],filter[4],mul_out[1735][23]);
mul_8x8bit m5207 (image[652],filter[5],mul_out[1735][24]);
mul_8x8bit m5208 (image[678],filter[6],mul_out[1736][22]);
mul_8x8bit m5209 (image[679],filter[7],mul_out[1736][23]);
mul_8x8bit m5210 (image[680],filter[8],mul_out[1736][24]);

adder_8bit ad578 (mul_out[1734][22],mul_out[1734][23],mul_out[1734][24],mul_out[1735][22],mul_out[1735][23],mul_out[1735][24],mul_out[1736][22],mul_out[1736][23],mul_out[1736][24],conv_out[578]);



mul_8x8bit m5211 (image[623],filter[0],mul_out[1737][22]);
mul_8x8bit m5212 (image[624],filter[1],mul_out[1737][23]);
mul_8x8bit m5213 (image[625],filter[2],mul_out[1737][24]);
mul_8x8bit m5214 (image[651],filter[3],mul_out[1738][22]);
mul_8x8bit m5215 (image[652],filter[4],mul_out[1738][23]);
mul_8x8bit m5216 (image[653],filter[5],mul_out[1738][24]);
mul_8x8bit m5217 (image[679],filter[6],mul_out[1739][22]);
mul_8x8bit m5218 (image[680],filter[7],mul_out[1739][23]);
mul_8x8bit m5219 (image[681],filter[8],mul_out[1739][24]);

adder_8bit ad579 (mul_out[1737][22],mul_out[1737][23],mul_out[1737][24],mul_out[1738][22],mul_out[1738][23],mul_out[1738][24],mul_out[1739][22],mul_out[1739][23],mul_out[1739][24],conv_out[579]);



mul_8x8bit m5220 (image[624],filter[0],mul_out[1740][22]);
mul_8x8bit m5221 (image[625],filter[1],mul_out[1740][23]);
mul_8x8bit m5222 (image[626],filter[2],mul_out[1740][24]);
mul_8x8bit m5223 (image[652],filter[3],mul_out[1741][22]);
mul_8x8bit m5224 (image[653],filter[4],mul_out[1741][23]);
mul_8x8bit m5225 (image[654],filter[5],mul_out[1741][24]);
mul_8x8bit m5226 (image[680],filter[6],mul_out[1742][22]);
mul_8x8bit m5227 (image[681],filter[7],mul_out[1742][23]);
mul_8x8bit m5228 (image[682],filter[8],mul_out[1742][24]);

adder_8bit ad580 (mul_out[1740][22],mul_out[1740][23],mul_out[1740][24],mul_out[1741][22],mul_out[1741][23],mul_out[1741][24],mul_out[1742][22],mul_out[1742][23],mul_out[1742][24],conv_out[580]);



mul_8x8bit m5229 (image[625],filter[0],mul_out[1743][22]);
mul_8x8bit m5230 (image[626],filter[1],mul_out[1743][23]);
mul_8x8bit m5231 (image[627],filter[2],mul_out[1743][24]);
mul_8x8bit m5232 (image[653],filter[3],mul_out[1744][22]);
mul_8x8bit m5233 (image[654],filter[4],mul_out[1744][23]);
mul_8x8bit m5234 (image[655],filter[5],mul_out[1744][24]);
mul_8x8bit m5235 (image[681],filter[6],mul_out[1745][22]);
mul_8x8bit m5236 (image[682],filter[7],mul_out[1745][23]);
mul_8x8bit m5237 (image[683],filter[8],mul_out[1745][24]);

adder_8bit ad581 (mul_out[1743][22],mul_out[1743][23],mul_out[1743][24],mul_out[1744][22],mul_out[1744][23],mul_out[1744][24],mul_out[1745][22],mul_out[1745][23],mul_out[1745][24],conv_out[581]);



mul_8x8bit m5238 (image[626],filter[0],mul_out[1746][22]);
mul_8x8bit m5239 (image[627],filter[1],mul_out[1746][23]);
mul_8x8bit m5240 (image[628],filter[2],mul_out[1746][24]);
mul_8x8bit m5241 (image[654],filter[3],mul_out[1747][22]);
mul_8x8bit m5242 (image[655],filter[4],mul_out[1747][23]);
mul_8x8bit m5243 (image[656],filter[5],mul_out[1747][24]);
mul_8x8bit m5244 (image[682],filter[6],mul_out[1748][22]);
mul_8x8bit m5245 (image[683],filter[7],mul_out[1748][23]);
mul_8x8bit m5246 (image[684],filter[8],mul_out[1748][24]);

adder_8bit ad582 (mul_out[1746][22],mul_out[1746][23],mul_out[1746][24],mul_out[1747][22],mul_out[1747][23],mul_out[1747][24],mul_out[1748][22],mul_out[1748][23],mul_out[1748][24],conv_out[582]);



mul_8x8bit m5247 (image[627],filter[0],mul_out[1749][22]);
mul_8x8bit m5248 (image[628],filter[1],mul_out[1749][23]);
mul_8x8bit m5249 (image[629],filter[2],mul_out[1749][24]);
mul_8x8bit m5250 (image[655],filter[3],mul_out[1750][22]);
mul_8x8bit m5251 (image[656],filter[4],mul_out[1750][23]);
mul_8x8bit m5252 (image[657],filter[5],mul_out[1750][24]);
mul_8x8bit m5253 (image[683],filter[6],mul_out[1751][22]);
mul_8x8bit m5254 (image[684],filter[7],mul_out[1751][23]);
mul_8x8bit m5255 (image[685],filter[8],mul_out[1751][24]);

adder_8bit ad583 (mul_out[1749][22],mul_out[1749][23],mul_out[1749][24],mul_out[1750][22],mul_out[1750][23],mul_out[1750][24],mul_out[1751][22],mul_out[1751][23],mul_out[1751][24],conv_out[583]);



mul_8x8bit m5256 (image[628],filter[0],mul_out[1752][22]);
mul_8x8bit m5257 (image[629],filter[1],mul_out[1752][23]);
mul_8x8bit m5258 (image[630],filter[2],mul_out[1752][24]);
mul_8x8bit m5259 (image[656],filter[3],mul_out[1753][22]);
mul_8x8bit m5260 (image[657],filter[4],mul_out[1753][23]);
mul_8x8bit m5261 (image[658],filter[5],mul_out[1753][24]);
mul_8x8bit m5262 (image[684],filter[6],mul_out[1754][22]);
mul_8x8bit m5263 (image[685],filter[7],mul_out[1754][23]);
mul_8x8bit m5264 (image[686],filter[8],mul_out[1754][24]);

adder_8bit ad584 (mul_out[1752][22],mul_out[1752][23],mul_out[1752][24],mul_out[1753][22],mul_out[1753][23],mul_out[1753][24],mul_out[1754][22],mul_out[1754][23],mul_out[1754][24],conv_out[584]);



mul_8x8bit m5265 (image[629],filter[0],mul_out[1755][22]);
mul_8x8bit m5266 (image[630],filter[1],mul_out[1755][23]);
mul_8x8bit m5267 (image[631],filter[2],mul_out[1755][24]);
mul_8x8bit m5268 (image[657],filter[3],mul_out[1756][22]);
mul_8x8bit m5269 (image[658],filter[4],mul_out[1756][23]);
mul_8x8bit m5270 (image[659],filter[5],mul_out[1756][24]);
mul_8x8bit m5271 (image[685],filter[6],mul_out[1757][22]);
mul_8x8bit m5272 (image[686],filter[7],mul_out[1757][23]);
mul_8x8bit m5273 (image[687],filter[8],mul_out[1757][24]);

adder_8bit ad585 (mul_out[1755][22],mul_out[1755][23],mul_out[1755][24],mul_out[1756][22],mul_out[1756][23],mul_out[1756][24],mul_out[1757][22],mul_out[1757][23],mul_out[1757][24],conv_out[585]);



mul_8x8bit m5274 (image[630],filter[0],mul_out[1758][22]);
mul_8x8bit m5275 (image[631],filter[1],mul_out[1758][23]);
mul_8x8bit m5276 (image[632],filter[2],mul_out[1758][24]);
mul_8x8bit m5277 (image[658],filter[3],mul_out[1759][22]);
mul_8x8bit m5278 (image[659],filter[4],mul_out[1759][23]);
mul_8x8bit m5279 (image[660],filter[5],mul_out[1759][24]);
mul_8x8bit m5280 (image[686],filter[6],mul_out[1760][22]);
mul_8x8bit m5281 (image[687],filter[7],mul_out[1760][23]);
mul_8x8bit m5282 (image[688],filter[8],mul_out[1760][24]);

adder_8bit ad586 (mul_out[1758][22],mul_out[1758][23],mul_out[1758][24],mul_out[1759][22],mul_out[1759][23],mul_out[1759][24],mul_out[1760][22],mul_out[1760][23],mul_out[1760][24],conv_out[586]);



mul_8x8bit m5283 (image[631],filter[0],mul_out[1761][22]);
mul_8x8bit m5284 (image[632],filter[1],mul_out[1761][23]);
mul_8x8bit m5285 (image[633],filter[2],mul_out[1761][24]);
mul_8x8bit m5286 (image[659],filter[3],mul_out[1762][22]);
mul_8x8bit m5287 (image[660],filter[4],mul_out[1762][23]);
mul_8x8bit m5288 (image[661],filter[5],mul_out[1762][24]);
mul_8x8bit m5289 (image[687],filter[6],mul_out[1763][22]);
mul_8x8bit m5290 (image[688],filter[7],mul_out[1763][23]);
mul_8x8bit m5291 (image[689],filter[8],mul_out[1763][24]);

adder_8bit ad587 (mul_out[1761][22],mul_out[1761][23],mul_out[1761][24],mul_out[1762][22],mul_out[1762][23],mul_out[1762][24],mul_out[1763][22],mul_out[1763][23],mul_out[1763][24],conv_out[587]);



mul_8x8bit m5292 (image[632],filter[0],mul_out[1764][22]);
mul_8x8bit m5293 (image[633],filter[1],mul_out[1764][23]);
mul_8x8bit m5294 (image[634],filter[2],mul_out[1764][24]);
mul_8x8bit m5295 (image[660],filter[3],mul_out[1765][22]);
mul_8x8bit m5296 (image[661],filter[4],mul_out[1765][23]);
mul_8x8bit m5297 (image[662],filter[5],mul_out[1765][24]);
mul_8x8bit m5298 (image[688],filter[6],mul_out[1766][22]);
mul_8x8bit m5299 (image[689],filter[7],mul_out[1766][23]);
mul_8x8bit m5300 (image[690],filter[8],mul_out[1766][24]);

adder_8bit ad588 (mul_out[1764][22],mul_out[1764][23],mul_out[1764][24],mul_out[1765][22],mul_out[1765][23],mul_out[1765][24],mul_out[1766][22],mul_out[1766][23],mul_out[1766][24],conv_out[588]);



mul_8x8bit m5301 (image[633],filter[0],mul_out[1767][22]);
mul_8x8bit m5302 (image[634],filter[1],mul_out[1767][23]);
mul_8x8bit m5303 (image[635],filter[2],mul_out[1767][24]);
mul_8x8bit m5304 (image[661],filter[3],mul_out[1768][22]);
mul_8x8bit m5305 (image[662],filter[4],mul_out[1768][23]);
mul_8x8bit m5306 (image[663],filter[5],mul_out[1768][24]);
mul_8x8bit m5307 (image[689],filter[6],mul_out[1769][22]);
mul_8x8bit m5308 (image[690],filter[7],mul_out[1769][23]);
mul_8x8bit m5309 (image[691],filter[8],mul_out[1769][24]);

adder_8bit ad589 (mul_out[1767][22],mul_out[1767][23],mul_out[1767][24],mul_out[1768][22],mul_out[1768][23],mul_out[1768][24],mul_out[1769][22],mul_out[1769][23],mul_out[1769][24],conv_out[589]);



mul_8x8bit m5310 (image[634],filter[0],mul_out[1770][22]);
mul_8x8bit m5311 (image[635],filter[1],mul_out[1770][23]);
mul_8x8bit m5312 (image[636],filter[2],mul_out[1770][24]);
mul_8x8bit m5313 (image[662],filter[3],mul_out[1771][22]);
mul_8x8bit m5314 (image[663],filter[4],mul_out[1771][23]);
mul_8x8bit m5315 (image[664],filter[5],mul_out[1771][24]);
mul_8x8bit m5316 (image[690],filter[6],mul_out[1772][22]);
mul_8x8bit m5317 (image[691],filter[7],mul_out[1772][23]);
mul_8x8bit m5318 (image[692],filter[8],mul_out[1772][24]);

adder_8bit ad590 (mul_out[1770][22],mul_out[1770][23],mul_out[1770][24],mul_out[1771][22],mul_out[1771][23],mul_out[1771][24],mul_out[1772][22],mul_out[1772][23],mul_out[1772][24],conv_out[590]);



mul_8x8bit m5319 (image[635],filter[0],mul_out[1773][22]);
mul_8x8bit m5320 (image[636],filter[1],mul_out[1773][23]);
mul_8x8bit m5321 (image[637],filter[2],mul_out[1773][24]);
mul_8x8bit m5322 (image[663],filter[3],mul_out[1774][22]);
mul_8x8bit m5323 (image[664],filter[4],mul_out[1774][23]);
mul_8x8bit m5324 (image[665],filter[5],mul_out[1774][24]);
mul_8x8bit m5325 (image[691],filter[6],mul_out[1775][22]);
mul_8x8bit m5326 (image[692],filter[7],mul_out[1775][23]);
mul_8x8bit m5327 (image[693],filter[8],mul_out[1775][24]);

adder_8bit ad591 (mul_out[1773][22],mul_out[1773][23],mul_out[1773][24],mul_out[1774][22],mul_out[1774][23],mul_out[1774][24],mul_out[1775][22],mul_out[1775][23],mul_out[1775][24],conv_out[591]);



mul_8x8bit m5328 (image[636],filter[0],mul_out[1776][22]);
mul_8x8bit m5329 (image[637],filter[1],mul_out[1776][23]);
mul_8x8bit m5330 (image[638],filter[2],mul_out[1776][24]);
mul_8x8bit m5331 (image[664],filter[3],mul_out[1777][22]);
mul_8x8bit m5332 (image[665],filter[4],mul_out[1777][23]);
mul_8x8bit m5333 (image[666],filter[5],mul_out[1777][24]);
mul_8x8bit m5334 (image[692],filter[6],mul_out[1778][22]);
mul_8x8bit m5335 (image[693],filter[7],mul_out[1778][23]);
mul_8x8bit m5336 (image[694],filter[8],mul_out[1778][24]);

adder_8bit ad592 (mul_out[1776][22],mul_out[1776][23],mul_out[1776][24],mul_out[1777][22],mul_out[1777][23],mul_out[1777][24],mul_out[1778][22],mul_out[1778][23],mul_out[1778][24],conv_out[592]);



mul_8x8bit m5337 (image[637],filter[0],mul_out[1779][22]);
mul_8x8bit m5338 (image[638],filter[1],mul_out[1779][23]);
mul_8x8bit m5339 (image[639],filter[2],mul_out[1779][24]);
mul_8x8bit m5340 (image[665],filter[3],mul_out[1780][22]);
mul_8x8bit m5341 (image[666],filter[4],mul_out[1780][23]);
mul_8x8bit m5342 (image[667],filter[5],mul_out[1780][24]);
mul_8x8bit m5343 (image[693],filter[6],mul_out[1781][22]);
mul_8x8bit m5344 (image[694],filter[7],mul_out[1781][23]);
mul_8x8bit m5345 (image[695],filter[8],mul_out[1781][24]);

adder_8bit ad593 (mul_out[1779][22],mul_out[1779][23],mul_out[1779][24],mul_out[1780][22],mul_out[1780][23],mul_out[1780][24],mul_out[1781][22],mul_out[1781][23],mul_out[1781][24],conv_out[593]);



mul_8x8bit m5346 (image[638],filter[0],mul_out[1782][22]);
mul_8x8bit m5347 (image[639],filter[1],mul_out[1782][23]);
mul_8x8bit m5348 (image[640],filter[2],mul_out[1782][24]);
mul_8x8bit m5349 (image[666],filter[3],mul_out[1783][22]);
mul_8x8bit m5350 (image[667],filter[4],mul_out[1783][23]);
mul_8x8bit m5351 (image[668],filter[5],mul_out[1783][24]);
mul_8x8bit m5352 (image[694],filter[6],mul_out[1784][22]);
mul_8x8bit m5353 (image[695],filter[7],mul_out[1784][23]);
mul_8x8bit m5354 (image[696],filter[8],mul_out[1784][24]);

adder_8bit ad594 (mul_out[1782][22],mul_out[1782][23],mul_out[1782][24],mul_out[1783][22],mul_out[1783][23],mul_out[1783][24],mul_out[1784][22],mul_out[1784][23],mul_out[1784][24],conv_out[594]);



mul_8x8bit m5355 (image[639],filter[0],mul_out[1785][22]);
mul_8x8bit m5356 (image[640],filter[1],mul_out[1785][23]);
mul_8x8bit m5357 (image[641],filter[2],mul_out[1785][24]);
mul_8x8bit m5358 (image[667],filter[3],mul_out[1786][22]);
mul_8x8bit m5359 (image[668],filter[4],mul_out[1786][23]);
mul_8x8bit m5360 (image[669],filter[5],mul_out[1786][24]);
mul_8x8bit m5361 (image[695],filter[6],mul_out[1787][22]);
mul_8x8bit m5362 (image[696],filter[7],mul_out[1787][23]);
mul_8x8bit m5363 (image[697],filter[8],mul_out[1787][24]);

adder_8bit ad595 (mul_out[1785][22],mul_out[1785][23],mul_out[1785][24],mul_out[1786][22],mul_out[1786][23],mul_out[1786][24],mul_out[1787][22],mul_out[1787][23],mul_out[1787][24],conv_out[595]);



mul_8x8bit m5364 (image[640],filter[0],mul_out[1788][22]);
mul_8x8bit m5365 (image[641],filter[1],mul_out[1788][23]);
mul_8x8bit m5366 (image[642],filter[2],mul_out[1788][24]);
mul_8x8bit m5367 (image[668],filter[3],mul_out[1789][22]);
mul_8x8bit m5368 (image[669],filter[4],mul_out[1789][23]);
mul_8x8bit m5369 (image[670],filter[5],mul_out[1789][24]);
mul_8x8bit m5370 (image[696],filter[6],mul_out[1790][22]);
mul_8x8bit m5371 (image[697],filter[7],mul_out[1790][23]);
mul_8x8bit m5372 (image[698],filter[8],mul_out[1790][24]);

adder_8bit ad596 (mul_out[1788][22],mul_out[1788][23],mul_out[1788][24],mul_out[1789][22],mul_out[1789][23],mul_out[1789][24],mul_out[1790][22],mul_out[1790][23],mul_out[1790][24],conv_out[596]);



mul_8x8bit m5373 (image[641],filter[0],mul_out[1791][22]);
mul_8x8bit m5374 (image[642],filter[1],mul_out[1791][23]);
mul_8x8bit m5375 (image[643],filter[2],mul_out[1791][24]);
mul_8x8bit m5376 (image[669],filter[3],mul_out[1792][22]);
mul_8x8bit m5377 (image[670],filter[4],mul_out[1792][23]);
mul_8x8bit m5378 (image[671],filter[5],mul_out[1792][24]);
mul_8x8bit m5379 (image[697],filter[6],mul_out[1793][22]);
mul_8x8bit m5380 (image[698],filter[7],mul_out[1793][23]);
mul_8x8bit m5381 (image[699],filter[8],mul_out[1793][24]);

adder_8bit ad597 (mul_out[1791][22],mul_out[1791][23],mul_out[1791][24],mul_out[1792][22],mul_out[1792][23],mul_out[1792][24],mul_out[1793][22],mul_out[1793][23],mul_out[1793][24],conv_out[597]);



mul_8x8bit m5382 (image[644],filter[0],mul_out[1794][23]);
mul_8x8bit m5383 (image[645],filter[1],mul_out[1794][24]);
mul_8x8bit m5384 (image[646],filter[2],mul_out[1794][25]);
mul_8x8bit m5385 (image[672],filter[3],mul_out[1795][23]);
mul_8x8bit m5386 (image[673],filter[4],mul_out[1795][24]);
mul_8x8bit m5387 (image[674],filter[5],mul_out[1795][25]);
mul_8x8bit m5388 (image[700],filter[6],mul_out[1796][23]);
mul_8x8bit m5389 (image[701],filter[7],mul_out[1796][24]);
mul_8x8bit m5390 (image[702],filter[8],mul_out[1796][25]);

adder_8bit ad598 (mul_out[1794][23],mul_out[1794][24],mul_out[1794][25],mul_out[1795][23],mul_out[1795][24],mul_out[1795][25],mul_out[1796][23],mul_out[1796][24],mul_out[1796][25],conv_out[598]);



mul_8x8bit m5391 (image[645],filter[0],mul_out[1797][23]);
mul_8x8bit m5392 (image[646],filter[1],mul_out[1797][24]);
mul_8x8bit m5393 (image[647],filter[2],mul_out[1797][25]);
mul_8x8bit m5394 (image[673],filter[3],mul_out[1798][23]);
mul_8x8bit m5395 (image[674],filter[4],mul_out[1798][24]);
mul_8x8bit m5396 (image[675],filter[5],mul_out[1798][25]);
mul_8x8bit m5397 (image[701],filter[6],mul_out[1799][23]);
mul_8x8bit m5398 (image[702],filter[7],mul_out[1799][24]);
mul_8x8bit m5399 (image[703],filter[8],mul_out[1799][25]);

adder_8bit ad599 (mul_out[1797][23],mul_out[1797][24],mul_out[1797][25],mul_out[1798][23],mul_out[1798][24],mul_out[1798][25],mul_out[1799][23],mul_out[1799][24],mul_out[1799][25],conv_out[599]);



mul_8x8bit m5400 (image[646],filter[0],mul_out[1800][23]);
mul_8x8bit m5401 (image[647],filter[1],mul_out[1800][24]);
mul_8x8bit m5402 (image[648],filter[2],mul_out[1800][25]);
mul_8x8bit m5403 (image[674],filter[3],mul_out[1801][23]);
mul_8x8bit m5404 (image[675],filter[4],mul_out[1801][24]);
mul_8x8bit m5405 (image[676],filter[5],mul_out[1801][25]);
mul_8x8bit m5406 (image[702],filter[6],mul_out[1802][23]);
mul_8x8bit m5407 (image[703],filter[7],mul_out[1802][24]);
mul_8x8bit m5408 (image[704],filter[8],mul_out[1802][25]);

adder_8bit ad600 (mul_out[1800][23],mul_out[1800][24],mul_out[1800][25],mul_out[1801][23],mul_out[1801][24],mul_out[1801][25],mul_out[1802][23],mul_out[1802][24],mul_out[1802][25],conv_out[600]);



mul_8x8bit m5409 (image[647],filter[0],mul_out[1803][23]);
mul_8x8bit m5410 (image[648],filter[1],mul_out[1803][24]);
mul_8x8bit m5411 (image[649],filter[2],mul_out[1803][25]);
mul_8x8bit m5412 (image[675],filter[3],mul_out[1804][23]);
mul_8x8bit m5413 (image[676],filter[4],mul_out[1804][24]);
mul_8x8bit m5414 (image[677],filter[5],mul_out[1804][25]);
mul_8x8bit m5415 (image[703],filter[6],mul_out[1805][23]);
mul_8x8bit m5416 (image[704],filter[7],mul_out[1805][24]);
mul_8x8bit m5417 (image[705],filter[8],mul_out[1805][25]);

adder_8bit ad601 (mul_out[1803][23],mul_out[1803][24],mul_out[1803][25],mul_out[1804][23],mul_out[1804][24],mul_out[1804][25],mul_out[1805][23],mul_out[1805][24],mul_out[1805][25],conv_out[601]);



mul_8x8bit m5418 (image[648],filter[0],mul_out[1806][23]);
mul_8x8bit m5419 (image[649],filter[1],mul_out[1806][24]);
mul_8x8bit m5420 (image[650],filter[2],mul_out[1806][25]);
mul_8x8bit m5421 (image[676],filter[3],mul_out[1807][23]);
mul_8x8bit m5422 (image[677],filter[4],mul_out[1807][24]);
mul_8x8bit m5423 (image[678],filter[5],mul_out[1807][25]);
mul_8x8bit m5424 (image[704],filter[6],mul_out[1808][23]);
mul_8x8bit m5425 (image[705],filter[7],mul_out[1808][24]);
mul_8x8bit m5426 (image[706],filter[8],mul_out[1808][25]);

adder_8bit ad602 (mul_out[1806][23],mul_out[1806][24],mul_out[1806][25],mul_out[1807][23],mul_out[1807][24],mul_out[1807][25],mul_out[1808][23],mul_out[1808][24],mul_out[1808][25],conv_out[602]);



mul_8x8bit m5427 (image[649],filter[0],mul_out[1809][23]);
mul_8x8bit m5428 (image[650],filter[1],mul_out[1809][24]);
mul_8x8bit m5429 (image[651],filter[2],mul_out[1809][25]);
mul_8x8bit m5430 (image[677],filter[3],mul_out[1810][23]);
mul_8x8bit m5431 (image[678],filter[4],mul_out[1810][24]);
mul_8x8bit m5432 (image[679],filter[5],mul_out[1810][25]);
mul_8x8bit m5433 (image[705],filter[6],mul_out[1811][23]);
mul_8x8bit m5434 (image[706],filter[7],mul_out[1811][24]);
mul_8x8bit m5435 (image[707],filter[8],mul_out[1811][25]);

adder_8bit ad603 (mul_out[1809][23],mul_out[1809][24],mul_out[1809][25],mul_out[1810][23],mul_out[1810][24],mul_out[1810][25],mul_out[1811][23],mul_out[1811][24],mul_out[1811][25],conv_out[603]);



mul_8x8bit m5436 (image[650],filter[0],mul_out[1812][23]);
mul_8x8bit m5437 (image[651],filter[1],mul_out[1812][24]);
mul_8x8bit m5438 (image[652],filter[2],mul_out[1812][25]);
mul_8x8bit m5439 (image[678],filter[3],mul_out[1813][23]);
mul_8x8bit m5440 (image[679],filter[4],mul_out[1813][24]);
mul_8x8bit m5441 (image[680],filter[5],mul_out[1813][25]);
mul_8x8bit m5442 (image[706],filter[6],mul_out[1814][23]);
mul_8x8bit m5443 (image[707],filter[7],mul_out[1814][24]);
mul_8x8bit m5444 (image[708],filter[8],mul_out[1814][25]);

adder_8bit ad604 (mul_out[1812][23],mul_out[1812][24],mul_out[1812][25],mul_out[1813][23],mul_out[1813][24],mul_out[1813][25],mul_out[1814][23],mul_out[1814][24],mul_out[1814][25],conv_out[604]);



mul_8x8bit m5445 (image[651],filter[0],mul_out[1815][23]);
mul_8x8bit m5446 (image[652],filter[1],mul_out[1815][24]);
mul_8x8bit m5447 (image[653],filter[2],mul_out[1815][25]);
mul_8x8bit m5448 (image[679],filter[3],mul_out[1816][23]);
mul_8x8bit m5449 (image[680],filter[4],mul_out[1816][24]);
mul_8x8bit m5450 (image[681],filter[5],mul_out[1816][25]);
mul_8x8bit m5451 (image[707],filter[6],mul_out[1817][23]);
mul_8x8bit m5452 (image[708],filter[7],mul_out[1817][24]);
mul_8x8bit m5453 (image[709],filter[8],mul_out[1817][25]);

adder_8bit ad605 (mul_out[1815][23],mul_out[1815][24],mul_out[1815][25],mul_out[1816][23],mul_out[1816][24],mul_out[1816][25],mul_out[1817][23],mul_out[1817][24],mul_out[1817][25],conv_out[605]);



mul_8x8bit m5454 (image[652],filter[0],mul_out[1818][23]);
mul_8x8bit m5455 (image[653],filter[1],mul_out[1818][24]);
mul_8x8bit m5456 (image[654],filter[2],mul_out[1818][25]);
mul_8x8bit m5457 (image[680],filter[3],mul_out[1819][23]);
mul_8x8bit m5458 (image[681],filter[4],mul_out[1819][24]);
mul_8x8bit m5459 (image[682],filter[5],mul_out[1819][25]);
mul_8x8bit m5460 (image[708],filter[6],mul_out[1820][23]);
mul_8x8bit m5461 (image[709],filter[7],mul_out[1820][24]);
mul_8x8bit m5462 (image[710],filter[8],mul_out[1820][25]);

adder_8bit ad606 (mul_out[1818][23],mul_out[1818][24],mul_out[1818][25],mul_out[1819][23],mul_out[1819][24],mul_out[1819][25],mul_out[1820][23],mul_out[1820][24],mul_out[1820][25],conv_out[606]);



mul_8x8bit m5463 (image[653],filter[0],mul_out[1821][23]);
mul_8x8bit m5464 (image[654],filter[1],mul_out[1821][24]);
mul_8x8bit m5465 (image[655],filter[2],mul_out[1821][25]);
mul_8x8bit m5466 (image[681],filter[3],mul_out[1822][23]);
mul_8x8bit m5467 (image[682],filter[4],mul_out[1822][24]);
mul_8x8bit m5468 (image[683],filter[5],mul_out[1822][25]);
mul_8x8bit m5469 (image[709],filter[6],mul_out[1823][23]);
mul_8x8bit m5470 (image[710],filter[7],mul_out[1823][24]);
mul_8x8bit m5471 (image[711],filter[8],mul_out[1823][25]);

adder_8bit ad607 (mul_out[1821][23],mul_out[1821][24],mul_out[1821][25],mul_out[1822][23],mul_out[1822][24],mul_out[1822][25],mul_out[1823][23],mul_out[1823][24],mul_out[1823][25],conv_out[607]);



mul_8x8bit m5472 (image[654],filter[0],mul_out[1824][23]);
mul_8x8bit m5473 (image[655],filter[1],mul_out[1824][24]);
mul_8x8bit m5474 (image[656],filter[2],mul_out[1824][25]);
mul_8x8bit m5475 (image[682],filter[3],mul_out[1825][23]);
mul_8x8bit m5476 (image[683],filter[4],mul_out[1825][24]);
mul_8x8bit m5477 (image[684],filter[5],mul_out[1825][25]);
mul_8x8bit m5478 (image[710],filter[6],mul_out[1826][23]);
mul_8x8bit m5479 (image[711],filter[7],mul_out[1826][24]);
mul_8x8bit m5480 (image[712],filter[8],mul_out[1826][25]);

adder_8bit ad608 (mul_out[1824][23],mul_out[1824][24],mul_out[1824][25],mul_out[1825][23],mul_out[1825][24],mul_out[1825][25],mul_out[1826][23],mul_out[1826][24],mul_out[1826][25],conv_out[608]);



mul_8x8bit m5481 (image[655],filter[0],mul_out[1827][23]);
mul_8x8bit m5482 (image[656],filter[1],mul_out[1827][24]);
mul_8x8bit m5483 (image[657],filter[2],mul_out[1827][25]);
mul_8x8bit m5484 (image[683],filter[3],mul_out[1828][23]);
mul_8x8bit m5485 (image[684],filter[4],mul_out[1828][24]);
mul_8x8bit m5486 (image[685],filter[5],mul_out[1828][25]);
mul_8x8bit m5487 (image[711],filter[6],mul_out[1829][23]);
mul_8x8bit m5488 (image[712],filter[7],mul_out[1829][24]);
mul_8x8bit m5489 (image[713],filter[8],mul_out[1829][25]);

adder_8bit ad609 (mul_out[1827][23],mul_out[1827][24],mul_out[1827][25],mul_out[1828][23],mul_out[1828][24],mul_out[1828][25],mul_out[1829][23],mul_out[1829][24],mul_out[1829][25],conv_out[609]);



mul_8x8bit m5490 (image[656],filter[0],mul_out[1830][23]);
mul_8x8bit m5491 (image[657],filter[1],mul_out[1830][24]);
mul_8x8bit m5492 (image[658],filter[2],mul_out[1830][25]);
mul_8x8bit m5493 (image[684],filter[3],mul_out[1831][23]);
mul_8x8bit m5494 (image[685],filter[4],mul_out[1831][24]);
mul_8x8bit m5495 (image[686],filter[5],mul_out[1831][25]);
mul_8x8bit m5496 (image[712],filter[6],mul_out[1832][23]);
mul_8x8bit m5497 (image[713],filter[7],mul_out[1832][24]);
mul_8x8bit m5498 (image[714],filter[8],mul_out[1832][25]);

adder_8bit ad610 (mul_out[1830][23],mul_out[1830][24],mul_out[1830][25],mul_out[1831][23],mul_out[1831][24],mul_out[1831][25],mul_out[1832][23],mul_out[1832][24],mul_out[1832][25],conv_out[610]);



mul_8x8bit m5499 (image[657],filter[0],mul_out[1833][23]);
mul_8x8bit m5500 (image[658],filter[1],mul_out[1833][24]);
mul_8x8bit m5501 (image[659],filter[2],mul_out[1833][25]);
mul_8x8bit m5502 (image[685],filter[3],mul_out[1834][23]);
mul_8x8bit m5503 (image[686],filter[4],mul_out[1834][24]);
mul_8x8bit m5504 (image[687],filter[5],mul_out[1834][25]);
mul_8x8bit m5505 (image[713],filter[6],mul_out[1835][23]);
mul_8x8bit m5506 (image[714],filter[7],mul_out[1835][24]);
mul_8x8bit m5507 (image[715],filter[8],mul_out[1835][25]);

adder_8bit ad611 (mul_out[1833][23],mul_out[1833][24],mul_out[1833][25],mul_out[1834][23],mul_out[1834][24],mul_out[1834][25],mul_out[1835][23],mul_out[1835][24],mul_out[1835][25],conv_out[611]);



mul_8x8bit m5508 (image[658],filter[0],mul_out[1836][23]);
mul_8x8bit m5509 (image[659],filter[1],mul_out[1836][24]);
mul_8x8bit m5510 (image[660],filter[2],mul_out[1836][25]);
mul_8x8bit m5511 (image[686],filter[3],mul_out[1837][23]);
mul_8x8bit m5512 (image[687],filter[4],mul_out[1837][24]);
mul_8x8bit m5513 (image[688],filter[5],mul_out[1837][25]);
mul_8x8bit m5514 (image[714],filter[6],mul_out[1838][23]);
mul_8x8bit m5515 (image[715],filter[7],mul_out[1838][24]);
mul_8x8bit m5516 (image[716],filter[8],mul_out[1838][25]);

adder_8bit ad612 (mul_out[1836][23],mul_out[1836][24],mul_out[1836][25],mul_out[1837][23],mul_out[1837][24],mul_out[1837][25],mul_out[1838][23],mul_out[1838][24],mul_out[1838][25],conv_out[612]);



mul_8x8bit m5517 (image[659],filter[0],mul_out[1839][23]);
mul_8x8bit m5518 (image[660],filter[1],mul_out[1839][24]);
mul_8x8bit m5519 (image[661],filter[2],mul_out[1839][25]);
mul_8x8bit m5520 (image[687],filter[3],mul_out[1840][23]);
mul_8x8bit m5521 (image[688],filter[4],mul_out[1840][24]);
mul_8x8bit m5522 (image[689],filter[5],mul_out[1840][25]);
mul_8x8bit m5523 (image[715],filter[6],mul_out[1841][23]);
mul_8x8bit m5524 (image[716],filter[7],mul_out[1841][24]);
mul_8x8bit m5525 (image[717],filter[8],mul_out[1841][25]);

adder_8bit ad613 (mul_out[1839][23],mul_out[1839][24],mul_out[1839][25],mul_out[1840][23],mul_out[1840][24],mul_out[1840][25],mul_out[1841][23],mul_out[1841][24],mul_out[1841][25],conv_out[613]);



mul_8x8bit m5526 (image[660],filter[0],mul_out[1842][23]);
mul_8x8bit m5527 (image[661],filter[1],mul_out[1842][24]);
mul_8x8bit m5528 (image[662],filter[2],mul_out[1842][25]);
mul_8x8bit m5529 (image[688],filter[3],mul_out[1843][23]);
mul_8x8bit m5530 (image[689],filter[4],mul_out[1843][24]);
mul_8x8bit m5531 (image[690],filter[5],mul_out[1843][25]);
mul_8x8bit m5532 (image[716],filter[6],mul_out[1844][23]);
mul_8x8bit m5533 (image[717],filter[7],mul_out[1844][24]);
mul_8x8bit m5534 (image[718],filter[8],mul_out[1844][25]);

adder_8bit ad614 (mul_out[1842][23],mul_out[1842][24],mul_out[1842][25],mul_out[1843][23],mul_out[1843][24],mul_out[1843][25],mul_out[1844][23],mul_out[1844][24],mul_out[1844][25],conv_out[614]);



mul_8x8bit m5535 (image[661],filter[0],mul_out[1845][23]);
mul_8x8bit m5536 (image[662],filter[1],mul_out[1845][24]);
mul_8x8bit m5537 (image[663],filter[2],mul_out[1845][25]);
mul_8x8bit m5538 (image[689],filter[3],mul_out[1846][23]);
mul_8x8bit m5539 (image[690],filter[4],mul_out[1846][24]);
mul_8x8bit m5540 (image[691],filter[5],mul_out[1846][25]);
mul_8x8bit m5541 (image[717],filter[6],mul_out[1847][23]);
mul_8x8bit m5542 (image[718],filter[7],mul_out[1847][24]);
mul_8x8bit m5543 (image[719],filter[8],mul_out[1847][25]);

adder_8bit ad615 (mul_out[1845][23],mul_out[1845][24],mul_out[1845][25],mul_out[1846][23],mul_out[1846][24],mul_out[1846][25],mul_out[1847][23],mul_out[1847][24],mul_out[1847][25],conv_out[615]);



mul_8x8bit m5544 (image[662],filter[0],mul_out[1848][23]);
mul_8x8bit m5545 (image[663],filter[1],mul_out[1848][24]);
mul_8x8bit m5546 (image[664],filter[2],mul_out[1848][25]);
mul_8x8bit m5547 (image[690],filter[3],mul_out[1849][23]);
mul_8x8bit m5548 (image[691],filter[4],mul_out[1849][24]);
mul_8x8bit m5549 (image[692],filter[5],mul_out[1849][25]);
mul_8x8bit m5550 (image[718],filter[6],mul_out[1850][23]);
mul_8x8bit m5551 (image[719],filter[7],mul_out[1850][24]);
mul_8x8bit m5552 (image[720],filter[8],mul_out[1850][25]);

adder_8bit ad616 (mul_out[1848][23],mul_out[1848][24],mul_out[1848][25],mul_out[1849][23],mul_out[1849][24],mul_out[1849][25],mul_out[1850][23],mul_out[1850][24],mul_out[1850][25],conv_out[616]);



mul_8x8bit m5553 (image[663],filter[0],mul_out[1851][23]);
mul_8x8bit m5554 (image[664],filter[1],mul_out[1851][24]);
mul_8x8bit m5555 (image[665],filter[2],mul_out[1851][25]);
mul_8x8bit m5556 (image[691],filter[3],mul_out[1852][23]);
mul_8x8bit m5557 (image[692],filter[4],mul_out[1852][24]);
mul_8x8bit m5558 (image[693],filter[5],mul_out[1852][25]);
mul_8x8bit m5559 (image[719],filter[6],mul_out[1853][23]);
mul_8x8bit m5560 (image[720],filter[7],mul_out[1853][24]);
mul_8x8bit m5561 (image[721],filter[8],mul_out[1853][25]);

adder_8bit ad617 (mul_out[1851][23],mul_out[1851][24],mul_out[1851][25],mul_out[1852][23],mul_out[1852][24],mul_out[1852][25],mul_out[1853][23],mul_out[1853][24],mul_out[1853][25],conv_out[617]);



mul_8x8bit m5562 (image[664],filter[0],mul_out[1854][23]);
mul_8x8bit m5563 (image[665],filter[1],mul_out[1854][24]);
mul_8x8bit m5564 (image[666],filter[2],mul_out[1854][25]);
mul_8x8bit m5565 (image[692],filter[3],mul_out[1855][23]);
mul_8x8bit m5566 (image[693],filter[4],mul_out[1855][24]);
mul_8x8bit m5567 (image[694],filter[5],mul_out[1855][25]);
mul_8x8bit m5568 (image[720],filter[6],mul_out[1856][23]);
mul_8x8bit m5569 (image[721],filter[7],mul_out[1856][24]);
mul_8x8bit m5570 (image[722],filter[8],mul_out[1856][25]);

adder_8bit ad618 (mul_out[1854][23],mul_out[1854][24],mul_out[1854][25],mul_out[1855][23],mul_out[1855][24],mul_out[1855][25],mul_out[1856][23],mul_out[1856][24],mul_out[1856][25],conv_out[618]);



mul_8x8bit m5571 (image[665],filter[0],mul_out[1857][23]);
mul_8x8bit m5572 (image[666],filter[1],mul_out[1857][24]);
mul_8x8bit m5573 (image[667],filter[2],mul_out[1857][25]);
mul_8x8bit m5574 (image[693],filter[3],mul_out[1858][23]);
mul_8x8bit m5575 (image[694],filter[4],mul_out[1858][24]);
mul_8x8bit m5576 (image[695],filter[5],mul_out[1858][25]);
mul_8x8bit m5577 (image[721],filter[6],mul_out[1859][23]);
mul_8x8bit m5578 (image[722],filter[7],mul_out[1859][24]);
mul_8x8bit m5579 (image[723],filter[8],mul_out[1859][25]);

adder_8bit ad619 (mul_out[1857][23],mul_out[1857][24],mul_out[1857][25],mul_out[1858][23],mul_out[1858][24],mul_out[1858][25],mul_out[1859][23],mul_out[1859][24],mul_out[1859][25],conv_out[619]);



mul_8x8bit m5580 (image[666],filter[0],mul_out[1860][23]);
mul_8x8bit m5581 (image[667],filter[1],mul_out[1860][24]);
mul_8x8bit m5582 (image[668],filter[2],mul_out[1860][25]);
mul_8x8bit m5583 (image[694],filter[3],mul_out[1861][23]);
mul_8x8bit m5584 (image[695],filter[4],mul_out[1861][24]);
mul_8x8bit m5585 (image[696],filter[5],mul_out[1861][25]);
mul_8x8bit m5586 (image[722],filter[6],mul_out[1862][23]);
mul_8x8bit m5587 (image[723],filter[7],mul_out[1862][24]);
mul_8x8bit m5588 (image[724],filter[8],mul_out[1862][25]);

adder_8bit ad620 (mul_out[1860][23],mul_out[1860][24],mul_out[1860][25],mul_out[1861][23],mul_out[1861][24],mul_out[1861][25],mul_out[1862][23],mul_out[1862][24],mul_out[1862][25],conv_out[620]);



mul_8x8bit m5589 (image[667],filter[0],mul_out[1863][23]);
mul_8x8bit m5590 (image[668],filter[1],mul_out[1863][24]);
mul_8x8bit m5591 (image[669],filter[2],mul_out[1863][25]);
mul_8x8bit m5592 (image[695],filter[3],mul_out[1864][23]);
mul_8x8bit m5593 (image[696],filter[4],mul_out[1864][24]);
mul_8x8bit m5594 (image[697],filter[5],mul_out[1864][25]);
mul_8x8bit m5595 (image[723],filter[6],mul_out[1865][23]);
mul_8x8bit m5596 (image[724],filter[7],mul_out[1865][24]);
mul_8x8bit m5597 (image[725],filter[8],mul_out[1865][25]);

adder_8bit ad621 (mul_out[1863][23],mul_out[1863][24],mul_out[1863][25],mul_out[1864][23],mul_out[1864][24],mul_out[1864][25],mul_out[1865][23],mul_out[1865][24],mul_out[1865][25],conv_out[621]);



mul_8x8bit m5598 (image[668],filter[0],mul_out[1866][23]);
mul_8x8bit m5599 (image[669],filter[1],mul_out[1866][24]);
mul_8x8bit m5600 (image[670],filter[2],mul_out[1866][25]);
mul_8x8bit m5601 (image[696],filter[3],mul_out[1867][23]);
mul_8x8bit m5602 (image[697],filter[4],mul_out[1867][24]);
mul_8x8bit m5603 (image[698],filter[5],mul_out[1867][25]);
mul_8x8bit m5604 (image[724],filter[6],mul_out[1868][23]);
mul_8x8bit m5605 (image[725],filter[7],mul_out[1868][24]);
mul_8x8bit m5606 (image[726],filter[8],mul_out[1868][25]);

adder_8bit ad622 (mul_out[1866][23],mul_out[1866][24],mul_out[1866][25],mul_out[1867][23],mul_out[1867][24],mul_out[1867][25],mul_out[1868][23],mul_out[1868][24],mul_out[1868][25],conv_out[622]);



mul_8x8bit m5607 (image[669],filter[0],mul_out[1869][23]);
mul_8x8bit m5608 (image[670],filter[1],mul_out[1869][24]);
mul_8x8bit m5609 (image[671],filter[2],mul_out[1869][25]);
mul_8x8bit m5610 (image[697],filter[3],mul_out[1870][23]);
mul_8x8bit m5611 (image[698],filter[4],mul_out[1870][24]);
mul_8x8bit m5612 (image[699],filter[5],mul_out[1870][25]);
mul_8x8bit m5613 (image[725],filter[6],mul_out[1871][23]);
mul_8x8bit m5614 (image[726],filter[7],mul_out[1871][24]);
mul_8x8bit m5615 (image[727],filter[8],mul_out[1871][25]);

adder_8bit ad623 (mul_out[1869][23],mul_out[1869][24],mul_out[1869][25],mul_out[1870][23],mul_out[1870][24],mul_out[1870][25],mul_out[1871][23],mul_out[1871][24],mul_out[1871][25],conv_out[623]);



mul_8x8bit m5616 (image[672],filter[0],mul_out[1872][24]);
mul_8x8bit m5617 (image[673],filter[1],mul_out[1872][25]);
mul_8x8bit m5618 (image[674],filter[2],mul_out[1872][26]);
mul_8x8bit m5619 (image[700],filter[3],mul_out[1873][24]);
mul_8x8bit m5620 (image[701],filter[4],mul_out[1873][25]);
mul_8x8bit m5621 (image[702],filter[5],mul_out[1873][26]);
mul_8x8bit m5622 (image[728],filter[6],mul_out[1874][24]);
mul_8x8bit m5623 (image[729],filter[7],mul_out[1874][25]);
mul_8x8bit m5624 (image[730],filter[8],mul_out[1874][26]);

adder_8bit ad624 (mul_out[1872][24],mul_out[1872][25],mul_out[1872][26],mul_out[1873][24],mul_out[1873][25],mul_out[1873][26],mul_out[1874][24],mul_out[1874][25],mul_out[1874][26],conv_out[624]);



mul_8x8bit m5625 (image[673],filter[0],mul_out[1875][24]);
mul_8x8bit m5626 (image[674],filter[1],mul_out[1875][25]);
mul_8x8bit m5627 (image[675],filter[2],mul_out[1875][26]);
mul_8x8bit m5628 (image[701],filter[3],mul_out[1876][24]);
mul_8x8bit m5629 (image[702],filter[4],mul_out[1876][25]);
mul_8x8bit m5630 (image[703],filter[5],mul_out[1876][26]);
mul_8x8bit m5631 (image[729],filter[6],mul_out[1877][24]);
mul_8x8bit m5632 (image[730],filter[7],mul_out[1877][25]);
mul_8x8bit m5633 (image[731],filter[8],mul_out[1877][26]);

adder_8bit ad625 (mul_out[1875][24],mul_out[1875][25],mul_out[1875][26],mul_out[1876][24],mul_out[1876][25],mul_out[1876][26],mul_out[1877][24],mul_out[1877][25],mul_out[1877][26],conv_out[625]);



mul_8x8bit m5634 (image[674],filter[0],mul_out[1878][24]);
mul_8x8bit m5635 (image[675],filter[1],mul_out[1878][25]);
mul_8x8bit m5636 (image[676],filter[2],mul_out[1878][26]);
mul_8x8bit m5637 (image[702],filter[3],mul_out[1879][24]);
mul_8x8bit m5638 (image[703],filter[4],mul_out[1879][25]);
mul_8x8bit m5639 (image[704],filter[5],mul_out[1879][26]);
mul_8x8bit m5640 (image[730],filter[6],mul_out[1880][24]);
mul_8x8bit m5641 (image[731],filter[7],mul_out[1880][25]);
mul_8x8bit m5642 (image[732],filter[8],mul_out[1880][26]);

adder_8bit ad626 (mul_out[1878][24],mul_out[1878][25],mul_out[1878][26],mul_out[1879][24],mul_out[1879][25],mul_out[1879][26],mul_out[1880][24],mul_out[1880][25],mul_out[1880][26],conv_out[626]);



mul_8x8bit m5643 (image[675],filter[0],mul_out[1881][24]);
mul_8x8bit m5644 (image[676],filter[1],mul_out[1881][25]);
mul_8x8bit m5645 (image[677],filter[2],mul_out[1881][26]);
mul_8x8bit m5646 (image[703],filter[3],mul_out[1882][24]);
mul_8x8bit m5647 (image[704],filter[4],mul_out[1882][25]);
mul_8x8bit m5648 (image[705],filter[5],mul_out[1882][26]);
mul_8x8bit m5649 (image[731],filter[6],mul_out[1883][24]);
mul_8x8bit m5650 (image[732],filter[7],mul_out[1883][25]);
mul_8x8bit m5651 (image[733],filter[8],mul_out[1883][26]);

adder_8bit ad627 (mul_out[1881][24],mul_out[1881][25],mul_out[1881][26],mul_out[1882][24],mul_out[1882][25],mul_out[1882][26],mul_out[1883][24],mul_out[1883][25],mul_out[1883][26],conv_out[627]);



mul_8x8bit m5652 (image[676],filter[0],mul_out[1884][24]);
mul_8x8bit m5653 (image[677],filter[1],mul_out[1884][25]);
mul_8x8bit m5654 (image[678],filter[2],mul_out[1884][26]);
mul_8x8bit m5655 (image[704],filter[3],mul_out[1885][24]);
mul_8x8bit m5656 (image[705],filter[4],mul_out[1885][25]);
mul_8x8bit m5657 (image[706],filter[5],mul_out[1885][26]);
mul_8x8bit m5658 (image[732],filter[6],mul_out[1886][24]);
mul_8x8bit m5659 (image[733],filter[7],mul_out[1886][25]);
mul_8x8bit m5660 (image[734],filter[8],mul_out[1886][26]);

adder_8bit ad628 (mul_out[1884][24],mul_out[1884][25],mul_out[1884][26],mul_out[1885][24],mul_out[1885][25],mul_out[1885][26],mul_out[1886][24],mul_out[1886][25],mul_out[1886][26],conv_out[628]);



mul_8x8bit m5661 (image[677],filter[0],mul_out[1887][24]);
mul_8x8bit m5662 (image[678],filter[1],mul_out[1887][25]);
mul_8x8bit m5663 (image[679],filter[2],mul_out[1887][26]);
mul_8x8bit m5664 (image[705],filter[3],mul_out[1888][24]);
mul_8x8bit m5665 (image[706],filter[4],mul_out[1888][25]);
mul_8x8bit m5666 (image[707],filter[5],mul_out[1888][26]);
mul_8x8bit m5667 (image[733],filter[6],mul_out[1889][24]);
mul_8x8bit m5668 (image[734],filter[7],mul_out[1889][25]);
mul_8x8bit m5669 (image[735],filter[8],mul_out[1889][26]);

adder_8bit ad629 (mul_out[1887][24],mul_out[1887][25],mul_out[1887][26],mul_out[1888][24],mul_out[1888][25],mul_out[1888][26],mul_out[1889][24],mul_out[1889][25],mul_out[1889][26],conv_out[629]);



mul_8x8bit m5670 (image[678],filter[0],mul_out[1890][24]);
mul_8x8bit m5671 (image[679],filter[1],mul_out[1890][25]);
mul_8x8bit m5672 (image[680],filter[2],mul_out[1890][26]);
mul_8x8bit m5673 (image[706],filter[3],mul_out[1891][24]);
mul_8x8bit m5674 (image[707],filter[4],mul_out[1891][25]);
mul_8x8bit m5675 (image[708],filter[5],mul_out[1891][26]);
mul_8x8bit m5676 (image[734],filter[6],mul_out[1892][24]);
mul_8x8bit m5677 (image[735],filter[7],mul_out[1892][25]);
mul_8x8bit m5678 (image[736],filter[8],mul_out[1892][26]);

adder_8bit ad630 (mul_out[1890][24],mul_out[1890][25],mul_out[1890][26],mul_out[1891][24],mul_out[1891][25],mul_out[1891][26],mul_out[1892][24],mul_out[1892][25],mul_out[1892][26],conv_out[630]);



mul_8x8bit m5679 (image[679],filter[0],mul_out[1893][24]);
mul_8x8bit m5680 (image[680],filter[1],mul_out[1893][25]);
mul_8x8bit m5681 (image[681],filter[2],mul_out[1893][26]);
mul_8x8bit m5682 (image[707],filter[3],mul_out[1894][24]);
mul_8x8bit m5683 (image[708],filter[4],mul_out[1894][25]);
mul_8x8bit m5684 (image[709],filter[5],mul_out[1894][26]);
mul_8x8bit m5685 (image[735],filter[6],mul_out[1895][24]);
mul_8x8bit m5686 (image[736],filter[7],mul_out[1895][25]);
mul_8x8bit m5687 (image[737],filter[8],mul_out[1895][26]);

adder_8bit ad631 (mul_out[1893][24],mul_out[1893][25],mul_out[1893][26],mul_out[1894][24],mul_out[1894][25],mul_out[1894][26],mul_out[1895][24],mul_out[1895][25],mul_out[1895][26],conv_out[631]);



mul_8x8bit m5688 (image[680],filter[0],mul_out[1896][24]);
mul_8x8bit m5689 (image[681],filter[1],mul_out[1896][25]);
mul_8x8bit m5690 (image[682],filter[2],mul_out[1896][26]);
mul_8x8bit m5691 (image[708],filter[3],mul_out[1897][24]);
mul_8x8bit m5692 (image[709],filter[4],mul_out[1897][25]);
mul_8x8bit m5693 (image[710],filter[5],mul_out[1897][26]);
mul_8x8bit m5694 (image[736],filter[6],mul_out[1898][24]);
mul_8x8bit m5695 (image[737],filter[7],mul_out[1898][25]);
mul_8x8bit m5696 (image[738],filter[8],mul_out[1898][26]);

adder_8bit ad632 (mul_out[1896][24],mul_out[1896][25],mul_out[1896][26],mul_out[1897][24],mul_out[1897][25],mul_out[1897][26],mul_out[1898][24],mul_out[1898][25],mul_out[1898][26],conv_out[632]);



mul_8x8bit m5697 (image[681],filter[0],mul_out[1899][24]);
mul_8x8bit m5698 (image[682],filter[1],mul_out[1899][25]);
mul_8x8bit m5699 (image[683],filter[2],mul_out[1899][26]);
mul_8x8bit m5700 (image[709],filter[3],mul_out[1900][24]);
mul_8x8bit m5701 (image[710],filter[4],mul_out[1900][25]);
mul_8x8bit m5702 (image[711],filter[5],mul_out[1900][26]);
mul_8x8bit m5703 (image[737],filter[6],mul_out[1901][24]);
mul_8x8bit m5704 (image[738],filter[7],mul_out[1901][25]);
mul_8x8bit m5705 (image[739],filter[8],mul_out[1901][26]);

adder_8bit ad633 (mul_out[1899][24],mul_out[1899][25],mul_out[1899][26],mul_out[1900][24],mul_out[1900][25],mul_out[1900][26],mul_out[1901][24],mul_out[1901][25],mul_out[1901][26],conv_out[633]);



mul_8x8bit m5706 (image[682],filter[0],mul_out[1902][24]);
mul_8x8bit m5707 (image[683],filter[1],mul_out[1902][25]);
mul_8x8bit m5708 (image[684],filter[2],mul_out[1902][26]);
mul_8x8bit m5709 (image[710],filter[3],mul_out[1903][24]);
mul_8x8bit m5710 (image[711],filter[4],mul_out[1903][25]);
mul_8x8bit m5711 (image[712],filter[5],mul_out[1903][26]);
mul_8x8bit m5712 (image[738],filter[6],mul_out[1904][24]);
mul_8x8bit m5713 (image[739],filter[7],mul_out[1904][25]);
mul_8x8bit m5714 (image[740],filter[8],mul_out[1904][26]);

adder_8bit ad634 (mul_out[1902][24],mul_out[1902][25],mul_out[1902][26],mul_out[1903][24],mul_out[1903][25],mul_out[1903][26],mul_out[1904][24],mul_out[1904][25],mul_out[1904][26],conv_out[634]);



mul_8x8bit m5715 (image[683],filter[0],mul_out[1905][24]);
mul_8x8bit m5716 (image[684],filter[1],mul_out[1905][25]);
mul_8x8bit m5717 (image[685],filter[2],mul_out[1905][26]);
mul_8x8bit m5718 (image[711],filter[3],mul_out[1906][24]);
mul_8x8bit m5719 (image[712],filter[4],mul_out[1906][25]);
mul_8x8bit m5720 (image[713],filter[5],mul_out[1906][26]);
mul_8x8bit m5721 (image[739],filter[6],mul_out[1907][24]);
mul_8x8bit m5722 (image[740],filter[7],mul_out[1907][25]);
mul_8x8bit m5723 (image[741],filter[8],mul_out[1907][26]);

adder_8bit ad635 (mul_out[1905][24],mul_out[1905][25],mul_out[1905][26],mul_out[1906][24],mul_out[1906][25],mul_out[1906][26],mul_out[1907][24],mul_out[1907][25],mul_out[1907][26],conv_out[635]);



mul_8x8bit m5724 (image[684],filter[0],mul_out[1908][24]);
mul_8x8bit m5725 (image[685],filter[1],mul_out[1908][25]);
mul_8x8bit m5726 (image[686],filter[2],mul_out[1908][26]);
mul_8x8bit m5727 (image[712],filter[3],mul_out[1909][24]);
mul_8x8bit m5728 (image[713],filter[4],mul_out[1909][25]);
mul_8x8bit m5729 (image[714],filter[5],mul_out[1909][26]);
mul_8x8bit m5730 (image[740],filter[6],mul_out[1910][24]);
mul_8x8bit m5731 (image[741],filter[7],mul_out[1910][25]);
mul_8x8bit m5732 (image[742],filter[8],mul_out[1910][26]);

adder_8bit ad636 (mul_out[1908][24],mul_out[1908][25],mul_out[1908][26],mul_out[1909][24],mul_out[1909][25],mul_out[1909][26],mul_out[1910][24],mul_out[1910][25],mul_out[1910][26],conv_out[636]);



mul_8x8bit m5733 (image[685],filter[0],mul_out[1911][24]);
mul_8x8bit m5734 (image[686],filter[1],mul_out[1911][25]);
mul_8x8bit m5735 (image[687],filter[2],mul_out[1911][26]);
mul_8x8bit m5736 (image[713],filter[3],mul_out[1912][24]);
mul_8x8bit m5737 (image[714],filter[4],mul_out[1912][25]);
mul_8x8bit m5738 (image[715],filter[5],mul_out[1912][26]);
mul_8x8bit m5739 (image[741],filter[6],mul_out[1913][24]);
mul_8x8bit m5740 (image[742],filter[7],mul_out[1913][25]);
mul_8x8bit m5741 (image[743],filter[8],mul_out[1913][26]);

adder_8bit ad637 (mul_out[1911][24],mul_out[1911][25],mul_out[1911][26],mul_out[1912][24],mul_out[1912][25],mul_out[1912][26],mul_out[1913][24],mul_out[1913][25],mul_out[1913][26],conv_out[637]);



mul_8x8bit m5742 (image[686],filter[0],mul_out[1914][24]);
mul_8x8bit m5743 (image[687],filter[1],mul_out[1914][25]);
mul_8x8bit m5744 (image[688],filter[2],mul_out[1914][26]);
mul_8x8bit m5745 (image[714],filter[3],mul_out[1915][24]);
mul_8x8bit m5746 (image[715],filter[4],mul_out[1915][25]);
mul_8x8bit m5747 (image[716],filter[5],mul_out[1915][26]);
mul_8x8bit m5748 (image[742],filter[6],mul_out[1916][24]);
mul_8x8bit m5749 (image[743],filter[7],mul_out[1916][25]);
mul_8x8bit m5750 (image[744],filter[8],mul_out[1916][26]);

adder_8bit ad638 (mul_out[1914][24],mul_out[1914][25],mul_out[1914][26],mul_out[1915][24],mul_out[1915][25],mul_out[1915][26],mul_out[1916][24],mul_out[1916][25],mul_out[1916][26],conv_out[638]);



mul_8x8bit m5751 (image[687],filter[0],mul_out[1917][24]);
mul_8x8bit m5752 (image[688],filter[1],mul_out[1917][25]);
mul_8x8bit m5753 (image[689],filter[2],mul_out[1917][26]);
mul_8x8bit m5754 (image[715],filter[3],mul_out[1918][24]);
mul_8x8bit m5755 (image[716],filter[4],mul_out[1918][25]);
mul_8x8bit m5756 (image[717],filter[5],mul_out[1918][26]);
mul_8x8bit m5757 (image[743],filter[6],mul_out[1919][24]);
mul_8x8bit m5758 (image[744],filter[7],mul_out[1919][25]);
mul_8x8bit m5759 (image[745],filter[8],mul_out[1919][26]);

adder_8bit ad639 (mul_out[1917][24],mul_out[1917][25],mul_out[1917][26],mul_out[1918][24],mul_out[1918][25],mul_out[1918][26],mul_out[1919][24],mul_out[1919][25],mul_out[1919][26],conv_out[639]);



mul_8x8bit m5760 (image[688],filter[0],mul_out[1920][24]);
mul_8x8bit m5761 (image[689],filter[1],mul_out[1920][25]);
mul_8x8bit m5762 (image[690],filter[2],mul_out[1920][26]);
mul_8x8bit m5763 (image[716],filter[3],mul_out[1921][24]);
mul_8x8bit m5764 (image[717],filter[4],mul_out[1921][25]);
mul_8x8bit m5765 (image[718],filter[5],mul_out[1921][26]);
mul_8x8bit m5766 (image[744],filter[6],mul_out[1922][24]);
mul_8x8bit m5767 (image[745],filter[7],mul_out[1922][25]);
mul_8x8bit m5768 (image[746],filter[8],mul_out[1922][26]);

adder_8bit ad640 (mul_out[1920][24],mul_out[1920][25],mul_out[1920][26],mul_out[1921][24],mul_out[1921][25],mul_out[1921][26],mul_out[1922][24],mul_out[1922][25],mul_out[1922][26],conv_out[640]);



mul_8x8bit m5769 (image[689],filter[0],mul_out[1923][24]);
mul_8x8bit m5770 (image[690],filter[1],mul_out[1923][25]);
mul_8x8bit m5771 (image[691],filter[2],mul_out[1923][26]);
mul_8x8bit m5772 (image[717],filter[3],mul_out[1924][24]);
mul_8x8bit m5773 (image[718],filter[4],mul_out[1924][25]);
mul_8x8bit m5774 (image[719],filter[5],mul_out[1924][26]);
mul_8x8bit m5775 (image[745],filter[6],mul_out[1925][24]);
mul_8x8bit m5776 (image[746],filter[7],mul_out[1925][25]);
mul_8x8bit m5777 (image[747],filter[8],mul_out[1925][26]);

adder_8bit ad641 (mul_out[1923][24],mul_out[1923][25],mul_out[1923][26],mul_out[1924][24],mul_out[1924][25],mul_out[1924][26],mul_out[1925][24],mul_out[1925][25],mul_out[1925][26],conv_out[641]);



mul_8x8bit m5778 (image[690],filter[0],mul_out[1926][24]);
mul_8x8bit m5779 (image[691],filter[1],mul_out[1926][25]);
mul_8x8bit m5780 (image[692],filter[2],mul_out[1926][26]);
mul_8x8bit m5781 (image[718],filter[3],mul_out[1927][24]);
mul_8x8bit m5782 (image[719],filter[4],mul_out[1927][25]);
mul_8x8bit m5783 (image[720],filter[5],mul_out[1927][26]);
mul_8x8bit m5784 (image[746],filter[6],mul_out[1928][24]);
mul_8x8bit m5785 (image[747],filter[7],mul_out[1928][25]);
mul_8x8bit m5786 (image[748],filter[8],mul_out[1928][26]);

adder_8bit ad642 (mul_out[1926][24],mul_out[1926][25],mul_out[1926][26],mul_out[1927][24],mul_out[1927][25],mul_out[1927][26],mul_out[1928][24],mul_out[1928][25],mul_out[1928][26],conv_out[642]);



mul_8x8bit m5787 (image[691],filter[0],mul_out[1929][24]);
mul_8x8bit m5788 (image[692],filter[1],mul_out[1929][25]);
mul_8x8bit m5789 (image[693],filter[2],mul_out[1929][26]);
mul_8x8bit m5790 (image[719],filter[3],mul_out[1930][24]);
mul_8x8bit m5791 (image[720],filter[4],mul_out[1930][25]);
mul_8x8bit m5792 (image[721],filter[5],mul_out[1930][26]);
mul_8x8bit m5793 (image[747],filter[6],mul_out[1931][24]);
mul_8x8bit m5794 (image[748],filter[7],mul_out[1931][25]);
mul_8x8bit m5795 (image[749],filter[8],mul_out[1931][26]);

adder_8bit ad643 (mul_out[1929][24],mul_out[1929][25],mul_out[1929][26],mul_out[1930][24],mul_out[1930][25],mul_out[1930][26],mul_out[1931][24],mul_out[1931][25],mul_out[1931][26],conv_out[643]);



mul_8x8bit m5796 (image[692],filter[0],mul_out[1932][24]);
mul_8x8bit m5797 (image[693],filter[1],mul_out[1932][25]);
mul_8x8bit m5798 (image[694],filter[2],mul_out[1932][26]);
mul_8x8bit m5799 (image[720],filter[3],mul_out[1933][24]);
mul_8x8bit m5800 (image[721],filter[4],mul_out[1933][25]);
mul_8x8bit m5801 (image[722],filter[5],mul_out[1933][26]);
mul_8x8bit m5802 (image[748],filter[6],mul_out[1934][24]);
mul_8x8bit m5803 (image[749],filter[7],mul_out[1934][25]);
mul_8x8bit m5804 (image[750],filter[8],mul_out[1934][26]);

adder_8bit ad644 (mul_out[1932][24],mul_out[1932][25],mul_out[1932][26],mul_out[1933][24],mul_out[1933][25],mul_out[1933][26],mul_out[1934][24],mul_out[1934][25],mul_out[1934][26],conv_out[644]);



mul_8x8bit m5805 (image[693],filter[0],mul_out[1935][24]);
mul_8x8bit m5806 (image[694],filter[1],mul_out[1935][25]);
mul_8x8bit m5807 (image[695],filter[2],mul_out[1935][26]);
mul_8x8bit m5808 (image[721],filter[3],mul_out[1936][24]);
mul_8x8bit m5809 (image[722],filter[4],mul_out[1936][25]);
mul_8x8bit m5810 (image[723],filter[5],mul_out[1936][26]);
mul_8x8bit m5811 (image[749],filter[6],mul_out[1937][24]);
mul_8x8bit m5812 (image[750],filter[7],mul_out[1937][25]);
mul_8x8bit m5813 (image[751],filter[8],mul_out[1937][26]);

adder_8bit ad645 (mul_out[1935][24],mul_out[1935][25],mul_out[1935][26],mul_out[1936][24],mul_out[1936][25],mul_out[1936][26],mul_out[1937][24],mul_out[1937][25],mul_out[1937][26],conv_out[645]);



mul_8x8bit m5814 (image[694],filter[0],mul_out[1938][24]);
mul_8x8bit m5815 (image[695],filter[1],mul_out[1938][25]);
mul_8x8bit m5816 (image[696],filter[2],mul_out[1938][26]);
mul_8x8bit m5817 (image[722],filter[3],mul_out[1939][24]);
mul_8x8bit m5818 (image[723],filter[4],mul_out[1939][25]);
mul_8x8bit m5819 (image[724],filter[5],mul_out[1939][26]);
mul_8x8bit m5820 (image[750],filter[6],mul_out[1940][24]);
mul_8x8bit m5821 (image[751],filter[7],mul_out[1940][25]);
mul_8x8bit m5822 (image[752],filter[8],mul_out[1940][26]);

adder_8bit ad646 (mul_out[1938][24],mul_out[1938][25],mul_out[1938][26],mul_out[1939][24],mul_out[1939][25],mul_out[1939][26],mul_out[1940][24],mul_out[1940][25],mul_out[1940][26],conv_out[646]);



mul_8x8bit m5823 (image[695],filter[0],mul_out[1941][24]);
mul_8x8bit m5824 (image[696],filter[1],mul_out[1941][25]);
mul_8x8bit m5825 (image[697],filter[2],mul_out[1941][26]);
mul_8x8bit m5826 (image[723],filter[3],mul_out[1942][24]);
mul_8x8bit m5827 (image[724],filter[4],mul_out[1942][25]);
mul_8x8bit m5828 (image[725],filter[5],mul_out[1942][26]);
mul_8x8bit m5829 (image[751],filter[6],mul_out[1943][24]);
mul_8x8bit m5830 (image[752],filter[7],mul_out[1943][25]);
mul_8x8bit m5831 (image[753],filter[8],mul_out[1943][26]);

adder_8bit ad647 (mul_out[1941][24],mul_out[1941][25],mul_out[1941][26],mul_out[1942][24],mul_out[1942][25],mul_out[1942][26],mul_out[1943][24],mul_out[1943][25],mul_out[1943][26],conv_out[647]);



mul_8x8bit m5832 (image[696],filter[0],mul_out[1944][24]);
mul_8x8bit m5833 (image[697],filter[1],mul_out[1944][25]);
mul_8x8bit m5834 (image[698],filter[2],mul_out[1944][26]);
mul_8x8bit m5835 (image[724],filter[3],mul_out[1945][24]);
mul_8x8bit m5836 (image[725],filter[4],mul_out[1945][25]);
mul_8x8bit m5837 (image[726],filter[5],mul_out[1945][26]);
mul_8x8bit m5838 (image[752],filter[6],mul_out[1946][24]);
mul_8x8bit m5839 (image[753],filter[7],mul_out[1946][25]);
mul_8x8bit m5840 (image[754],filter[8],mul_out[1946][26]);

adder_8bit ad648 (mul_out[1944][24],mul_out[1944][25],mul_out[1944][26],mul_out[1945][24],mul_out[1945][25],mul_out[1945][26],mul_out[1946][24],mul_out[1946][25],mul_out[1946][26],conv_out[648]);



mul_8x8bit m5841 (image[697],filter[0],mul_out[1947][24]);
mul_8x8bit m5842 (image[698],filter[1],mul_out[1947][25]);
mul_8x8bit m5843 (image[699],filter[2],mul_out[1947][26]);
mul_8x8bit m5844 (image[725],filter[3],mul_out[1948][24]);
mul_8x8bit m5845 (image[726],filter[4],mul_out[1948][25]);
mul_8x8bit m5846 (image[727],filter[5],mul_out[1948][26]);
mul_8x8bit m5847 (image[753],filter[6],mul_out[1949][24]);
mul_8x8bit m5848 (image[754],filter[7],mul_out[1949][25]);
mul_8x8bit m5849 (image[755],filter[8],mul_out[1949][26]);

adder_8bit ad649 (mul_out[1947][24],mul_out[1947][25],mul_out[1947][26],mul_out[1948][24],mul_out[1948][25],mul_out[1948][26],mul_out[1949][24],mul_out[1949][25],mul_out[1949][26],conv_out[649]);



mul_8x8bit m5850 (image[700],filter[0],mul_out[1950][25]);
mul_8x8bit m5851 (image[701],filter[1],mul_out[1950][26]);
mul_8x8bit m5852 (image[702],filter[2],mul_out[1950][27]);
mul_8x8bit m5853 (image[728],filter[3],mul_out[1951][25]);
mul_8x8bit m5854 (image[729],filter[4],mul_out[1951][26]);
mul_8x8bit m5855 (image[730],filter[5],mul_out[1951][27]);
mul_8x8bit m5856 (image[756],filter[6],mul_out[1952][25]);
mul_8x8bit m5857 (image[757],filter[7],mul_out[1952][26]);
mul_8x8bit m5858 (image[758],filter[8],mul_out[1952][27]);

adder_8bit ad650 (mul_out[1950][25],mul_out[1950][26],mul_out[1950][27],mul_out[1951][25],mul_out[1951][26],mul_out[1951][27],mul_out[1952][25],mul_out[1952][26],mul_out[1952][27],conv_out[650]);



mul_8x8bit m5859 (image[701],filter[0],mul_out[1953][25]);
mul_8x8bit m5860 (image[702],filter[1],mul_out[1953][26]);
mul_8x8bit m5861 (image[703],filter[2],mul_out[1953][27]);
mul_8x8bit m5862 (image[729],filter[3],mul_out[1954][25]);
mul_8x8bit m5863 (image[730],filter[4],mul_out[1954][26]);
mul_8x8bit m5864 (image[731],filter[5],mul_out[1954][27]);
mul_8x8bit m5865 (image[757],filter[6],mul_out[1955][25]);
mul_8x8bit m5866 (image[758],filter[7],mul_out[1955][26]);
mul_8x8bit m5867 (image[759],filter[8],mul_out[1955][27]);

adder_8bit ad651 (mul_out[1953][25],mul_out[1953][26],mul_out[1953][27],mul_out[1954][25],mul_out[1954][26],mul_out[1954][27],mul_out[1955][25],mul_out[1955][26],mul_out[1955][27],conv_out[651]);



mul_8x8bit m5868 (image[702],filter[0],mul_out[1956][25]);
mul_8x8bit m5869 (image[703],filter[1],mul_out[1956][26]);
mul_8x8bit m5870 (image[704],filter[2],mul_out[1956][27]);
mul_8x8bit m5871 (image[730],filter[3],mul_out[1957][25]);
mul_8x8bit m5872 (image[731],filter[4],mul_out[1957][26]);
mul_8x8bit m5873 (image[732],filter[5],mul_out[1957][27]);
mul_8x8bit m5874 (image[758],filter[6],mul_out[1958][25]);
mul_8x8bit m5875 (image[759],filter[7],mul_out[1958][26]);
mul_8x8bit m5876 (image[760],filter[8],mul_out[1958][27]);

adder_8bit ad652 (mul_out[1956][25],mul_out[1956][26],mul_out[1956][27],mul_out[1957][25],mul_out[1957][26],mul_out[1957][27],mul_out[1958][25],mul_out[1958][26],mul_out[1958][27],conv_out[652]);



mul_8x8bit m5877 (image[703],filter[0],mul_out[1959][25]);
mul_8x8bit m5878 (image[704],filter[1],mul_out[1959][26]);
mul_8x8bit m5879 (image[705],filter[2],mul_out[1959][27]);
mul_8x8bit m5880 (image[731],filter[3],mul_out[1960][25]);
mul_8x8bit m5881 (image[732],filter[4],mul_out[1960][26]);
mul_8x8bit m5882 (image[733],filter[5],mul_out[1960][27]);
mul_8x8bit m5883 (image[759],filter[6],mul_out[1961][25]);
mul_8x8bit m5884 (image[760],filter[7],mul_out[1961][26]);
mul_8x8bit m5885 (image[761],filter[8],mul_out[1961][27]);

adder_8bit ad653 (mul_out[1959][25],mul_out[1959][26],mul_out[1959][27],mul_out[1960][25],mul_out[1960][26],mul_out[1960][27],mul_out[1961][25],mul_out[1961][26],mul_out[1961][27],conv_out[653]);



mul_8x8bit m5886 (image[704],filter[0],mul_out[1962][25]);
mul_8x8bit m5887 (image[705],filter[1],mul_out[1962][26]);
mul_8x8bit m5888 (image[706],filter[2],mul_out[1962][27]);
mul_8x8bit m5889 (image[732],filter[3],mul_out[1963][25]);
mul_8x8bit m5890 (image[733],filter[4],mul_out[1963][26]);
mul_8x8bit m5891 (image[734],filter[5],mul_out[1963][27]);
mul_8x8bit m5892 (image[760],filter[6],mul_out[1964][25]);
mul_8x8bit m5893 (image[761],filter[7],mul_out[1964][26]);
mul_8x8bit m5894 (image[762],filter[8],mul_out[1964][27]);

adder_8bit ad654 (mul_out[1962][25],mul_out[1962][26],mul_out[1962][27],mul_out[1963][25],mul_out[1963][26],mul_out[1963][27],mul_out[1964][25],mul_out[1964][26],mul_out[1964][27],conv_out[654]);



mul_8x8bit m5895 (image[705],filter[0],mul_out[1965][25]);
mul_8x8bit m5896 (image[706],filter[1],mul_out[1965][26]);
mul_8x8bit m5897 (image[707],filter[2],mul_out[1965][27]);
mul_8x8bit m5898 (image[733],filter[3],mul_out[1966][25]);
mul_8x8bit m5899 (image[734],filter[4],mul_out[1966][26]);
mul_8x8bit m5900 (image[735],filter[5],mul_out[1966][27]);
mul_8x8bit m5901 (image[761],filter[6],mul_out[1967][25]);
mul_8x8bit m5902 (image[762],filter[7],mul_out[1967][26]);
mul_8x8bit m5903 (image[763],filter[8],mul_out[1967][27]);

adder_8bit ad655 (mul_out[1965][25],mul_out[1965][26],mul_out[1965][27],mul_out[1966][25],mul_out[1966][26],mul_out[1966][27],mul_out[1967][25],mul_out[1967][26],mul_out[1967][27],conv_out[655]);



mul_8x8bit m5904 (image[706],filter[0],mul_out[1968][25]);
mul_8x8bit m5905 (image[707],filter[1],mul_out[1968][26]);
mul_8x8bit m5906 (image[708],filter[2],mul_out[1968][27]);
mul_8x8bit m5907 (image[734],filter[3],mul_out[1969][25]);
mul_8x8bit m5908 (image[735],filter[4],mul_out[1969][26]);
mul_8x8bit m5909 (image[736],filter[5],mul_out[1969][27]);
mul_8x8bit m5910 (image[762],filter[6],mul_out[1970][25]);
mul_8x8bit m5911 (image[763],filter[7],mul_out[1970][26]);
mul_8x8bit m5912 (image[764],filter[8],mul_out[1970][27]);

adder_8bit ad656 (mul_out[1968][25],mul_out[1968][26],mul_out[1968][27],mul_out[1969][25],mul_out[1969][26],mul_out[1969][27],mul_out[1970][25],mul_out[1970][26],mul_out[1970][27],conv_out[656]);



mul_8x8bit m5913 (image[707],filter[0],mul_out[1971][25]);
mul_8x8bit m5914 (image[708],filter[1],mul_out[1971][26]);
mul_8x8bit m5915 (image[709],filter[2],mul_out[1971][27]);
mul_8x8bit m5916 (image[735],filter[3],mul_out[1972][25]);
mul_8x8bit m5917 (image[736],filter[4],mul_out[1972][26]);
mul_8x8bit m5918 (image[737],filter[5],mul_out[1972][27]);
mul_8x8bit m5919 (image[763],filter[6],mul_out[1973][25]);
mul_8x8bit m5920 (image[764],filter[7],mul_out[1973][26]);
mul_8x8bit m5921 (image[765],filter[8],mul_out[1973][27]);

adder_8bit ad657 (mul_out[1971][25],mul_out[1971][26],mul_out[1971][27],mul_out[1972][25],mul_out[1972][26],mul_out[1972][27],mul_out[1973][25],mul_out[1973][26],mul_out[1973][27],conv_out[657]);



mul_8x8bit m5922 (image[708],filter[0],mul_out[1974][25]);
mul_8x8bit m5923 (image[709],filter[1],mul_out[1974][26]);
mul_8x8bit m5924 (image[710],filter[2],mul_out[1974][27]);
mul_8x8bit m5925 (image[736],filter[3],mul_out[1975][25]);
mul_8x8bit m5926 (image[737],filter[4],mul_out[1975][26]);
mul_8x8bit m5927 (image[738],filter[5],mul_out[1975][27]);
mul_8x8bit m5928 (image[764],filter[6],mul_out[1976][25]);
mul_8x8bit m5929 (image[765],filter[7],mul_out[1976][26]);
mul_8x8bit m5930 (image[766],filter[8],mul_out[1976][27]);

adder_8bit ad658 (mul_out[1974][25],mul_out[1974][26],mul_out[1974][27],mul_out[1975][25],mul_out[1975][26],mul_out[1975][27],mul_out[1976][25],mul_out[1976][26],mul_out[1976][27],conv_out[658]);



mul_8x8bit m5931 (image[709],filter[0],mul_out[1977][25]);
mul_8x8bit m5932 (image[710],filter[1],mul_out[1977][26]);
mul_8x8bit m5933 (image[711],filter[2],mul_out[1977][27]);
mul_8x8bit m5934 (image[737],filter[3],mul_out[1978][25]);
mul_8x8bit m5935 (image[738],filter[4],mul_out[1978][26]);
mul_8x8bit m5936 (image[739],filter[5],mul_out[1978][27]);
mul_8x8bit m5937 (image[765],filter[6],mul_out[1979][25]);
mul_8x8bit m5938 (image[766],filter[7],mul_out[1979][26]);
mul_8x8bit m5939 (image[767],filter[8],mul_out[1979][27]);

adder_8bit ad659 (mul_out[1977][25],mul_out[1977][26],mul_out[1977][27],mul_out[1978][25],mul_out[1978][26],mul_out[1978][27],mul_out[1979][25],mul_out[1979][26],mul_out[1979][27],conv_out[659]);



mul_8x8bit m5940 (image[710],filter[0],mul_out[1980][25]);
mul_8x8bit m5941 (image[711],filter[1],mul_out[1980][26]);
mul_8x8bit m5942 (image[712],filter[2],mul_out[1980][27]);
mul_8x8bit m5943 (image[738],filter[3],mul_out[1981][25]);
mul_8x8bit m5944 (image[739],filter[4],mul_out[1981][26]);
mul_8x8bit m5945 (image[740],filter[5],mul_out[1981][27]);
mul_8x8bit m5946 (image[766],filter[6],mul_out[1982][25]);
mul_8x8bit m5947 (image[767],filter[7],mul_out[1982][26]);
mul_8x8bit m5948 (image[768],filter[8],mul_out[1982][27]);

adder_8bit ad660 (mul_out[1980][25],mul_out[1980][26],mul_out[1980][27],mul_out[1981][25],mul_out[1981][26],mul_out[1981][27],mul_out[1982][25],mul_out[1982][26],mul_out[1982][27],conv_out[660]);



mul_8x8bit m5949 (image[711],filter[0],mul_out[1983][25]);
mul_8x8bit m5950 (image[712],filter[1],mul_out[1983][26]);
mul_8x8bit m5951 (image[713],filter[2],mul_out[1983][27]);
mul_8x8bit m5952 (image[739],filter[3],mul_out[1984][25]);
mul_8x8bit m5953 (image[740],filter[4],mul_out[1984][26]);
mul_8x8bit m5954 (image[741],filter[5],mul_out[1984][27]);
mul_8x8bit m5955 (image[767],filter[6],mul_out[1985][25]);
mul_8x8bit m5956 (image[768],filter[7],mul_out[1985][26]);
mul_8x8bit m5957 (image[769],filter[8],mul_out[1985][27]);

adder_8bit ad661 (mul_out[1983][25],mul_out[1983][26],mul_out[1983][27],mul_out[1984][25],mul_out[1984][26],mul_out[1984][27],mul_out[1985][25],mul_out[1985][26],mul_out[1985][27],conv_out[661]);



mul_8x8bit m5958 (image[712],filter[0],mul_out[1986][25]);
mul_8x8bit m5959 (image[713],filter[1],mul_out[1986][26]);
mul_8x8bit m5960 (image[714],filter[2],mul_out[1986][27]);
mul_8x8bit m5961 (image[740],filter[3],mul_out[1987][25]);
mul_8x8bit m5962 (image[741],filter[4],mul_out[1987][26]);
mul_8x8bit m5963 (image[742],filter[5],mul_out[1987][27]);
mul_8x8bit m5964 (image[768],filter[6],mul_out[1988][25]);
mul_8x8bit m5965 (image[769],filter[7],mul_out[1988][26]);
mul_8x8bit m5966 (image[770],filter[8],mul_out[1988][27]);

adder_8bit ad662 (mul_out[1986][25],mul_out[1986][26],mul_out[1986][27],mul_out[1987][25],mul_out[1987][26],mul_out[1987][27],mul_out[1988][25],mul_out[1988][26],mul_out[1988][27],conv_out[662]);



mul_8x8bit m5967 (image[713],filter[0],mul_out[1989][25]);
mul_8x8bit m5968 (image[714],filter[1],mul_out[1989][26]);
mul_8x8bit m5969 (image[715],filter[2],mul_out[1989][27]);
mul_8x8bit m5970 (image[741],filter[3],mul_out[1990][25]);
mul_8x8bit m5971 (image[742],filter[4],mul_out[1990][26]);
mul_8x8bit m5972 (image[743],filter[5],mul_out[1990][27]);
mul_8x8bit m5973 (image[769],filter[6],mul_out[1991][25]);
mul_8x8bit m5974 (image[770],filter[7],mul_out[1991][26]);
mul_8x8bit m5975 (image[771],filter[8],mul_out[1991][27]);

adder_8bit ad663 (mul_out[1989][25],mul_out[1989][26],mul_out[1989][27],mul_out[1990][25],mul_out[1990][26],mul_out[1990][27],mul_out[1991][25],mul_out[1991][26],mul_out[1991][27],conv_out[663]);



mul_8x8bit m5976 (image[714],filter[0],mul_out[1992][25]);
mul_8x8bit m5977 (image[715],filter[1],mul_out[1992][26]);
mul_8x8bit m5978 (image[716],filter[2],mul_out[1992][27]);
mul_8x8bit m5979 (image[742],filter[3],mul_out[1993][25]);
mul_8x8bit m5980 (image[743],filter[4],mul_out[1993][26]);
mul_8x8bit m5981 (image[744],filter[5],mul_out[1993][27]);
mul_8x8bit m5982 (image[770],filter[6],mul_out[1994][25]);
mul_8x8bit m5983 (image[771],filter[7],mul_out[1994][26]);
mul_8x8bit m5984 (image[772],filter[8],mul_out[1994][27]);

adder_8bit ad664 (mul_out[1992][25],mul_out[1992][26],mul_out[1992][27],mul_out[1993][25],mul_out[1993][26],mul_out[1993][27],mul_out[1994][25],mul_out[1994][26],mul_out[1994][27],conv_out[664]);



mul_8x8bit m5985 (image[715],filter[0],mul_out[1995][25]);
mul_8x8bit m5986 (image[716],filter[1],mul_out[1995][26]);
mul_8x8bit m5987 (image[717],filter[2],mul_out[1995][27]);
mul_8x8bit m5988 (image[743],filter[3],mul_out[1996][25]);
mul_8x8bit m5989 (image[744],filter[4],mul_out[1996][26]);
mul_8x8bit m5990 (image[745],filter[5],mul_out[1996][27]);
mul_8x8bit m5991 (image[771],filter[6],mul_out[1997][25]);
mul_8x8bit m5992 (image[772],filter[7],mul_out[1997][26]);
mul_8x8bit m5993 (image[773],filter[8],mul_out[1997][27]);

adder_8bit ad665 (mul_out[1995][25],mul_out[1995][26],mul_out[1995][27],mul_out[1996][25],mul_out[1996][26],mul_out[1996][27],mul_out[1997][25],mul_out[1997][26],mul_out[1997][27],conv_out[665]);



mul_8x8bit m5994 (image[716],filter[0],mul_out[1998][25]);
mul_8x8bit m5995 (image[717],filter[1],mul_out[1998][26]);
mul_8x8bit m5996 (image[718],filter[2],mul_out[1998][27]);
mul_8x8bit m5997 (image[744],filter[3],mul_out[1999][25]);
mul_8x8bit m5998 (image[745],filter[4],mul_out[1999][26]);
mul_8x8bit m5999 (image[746],filter[5],mul_out[1999][27]);
mul_8x8bit m6000 (image[772],filter[6],mul_out[2000][25]);
mul_8x8bit m6001 (image[773],filter[7],mul_out[2000][26]);
mul_8x8bit m6002 (image[774],filter[8],mul_out[2000][27]);

adder_8bit ad666 (mul_out[1998][25],mul_out[1998][26],mul_out[1998][27],mul_out[1999][25],mul_out[1999][26],mul_out[1999][27],mul_out[2000][25],mul_out[2000][26],mul_out[2000][27],conv_out[666]);



mul_8x8bit m6003 (image[717],filter[0],mul_out[2001][25]);
mul_8x8bit m6004 (image[718],filter[1],mul_out[2001][26]);
mul_8x8bit m6005 (image[719],filter[2],mul_out[2001][27]);
mul_8x8bit m6006 (image[745],filter[3],mul_out[2002][25]);
mul_8x8bit m6007 (image[746],filter[4],mul_out[2002][26]);
mul_8x8bit m6008 (image[747],filter[5],mul_out[2002][27]);
mul_8x8bit m6009 (image[773],filter[6],mul_out[2003][25]);
mul_8x8bit m6010 (image[774],filter[7],mul_out[2003][26]);
mul_8x8bit m6011 (image[775],filter[8],mul_out[2003][27]);

adder_8bit ad667 (mul_out[2001][25],mul_out[2001][26],mul_out[2001][27],mul_out[2002][25],mul_out[2002][26],mul_out[2002][27],mul_out[2003][25],mul_out[2003][26],mul_out[2003][27],conv_out[667]);



mul_8x8bit m6012 (image[718],filter[0],mul_out[2004][25]);
mul_8x8bit m6013 (image[719],filter[1],mul_out[2004][26]);
mul_8x8bit m6014 (image[720],filter[2],mul_out[2004][27]);
mul_8x8bit m6015 (image[746],filter[3],mul_out[2005][25]);
mul_8x8bit m6016 (image[747],filter[4],mul_out[2005][26]);
mul_8x8bit m6017 (image[748],filter[5],mul_out[2005][27]);
mul_8x8bit m6018 (image[774],filter[6],mul_out[2006][25]);
mul_8x8bit m6019 (image[775],filter[7],mul_out[2006][26]);
mul_8x8bit m6020 (image[776],filter[8],mul_out[2006][27]);

adder_8bit ad668 (mul_out[2004][25],mul_out[2004][26],mul_out[2004][27],mul_out[2005][25],mul_out[2005][26],mul_out[2005][27],mul_out[2006][25],mul_out[2006][26],mul_out[2006][27],conv_out[668]);



mul_8x8bit m6021 (image[719],filter[0],mul_out[2007][25]);
mul_8x8bit m6022 (image[720],filter[1],mul_out[2007][26]);
mul_8x8bit m6023 (image[721],filter[2],mul_out[2007][27]);
mul_8x8bit m6024 (image[747],filter[3],mul_out[2008][25]);
mul_8x8bit m6025 (image[748],filter[4],mul_out[2008][26]);
mul_8x8bit m6026 (image[749],filter[5],mul_out[2008][27]);
mul_8x8bit m6027 (image[775],filter[6],mul_out[2009][25]);
mul_8x8bit m6028 (image[776],filter[7],mul_out[2009][26]);
mul_8x8bit m6029 (image[777],filter[8],mul_out[2009][27]);

adder_8bit ad669 (mul_out[2007][25],mul_out[2007][26],mul_out[2007][27],mul_out[2008][25],mul_out[2008][26],mul_out[2008][27],mul_out[2009][25],mul_out[2009][26],mul_out[2009][27],conv_out[669]);



mul_8x8bit m6030 (image[720],filter[0],mul_out[2010][25]);
mul_8x8bit m6031 (image[721],filter[1],mul_out[2010][26]);
mul_8x8bit m6032 (image[722],filter[2],mul_out[2010][27]);
mul_8x8bit m6033 (image[748],filter[3],mul_out[2011][25]);
mul_8x8bit m6034 (image[749],filter[4],mul_out[2011][26]);
mul_8x8bit m6035 (image[750],filter[5],mul_out[2011][27]);
mul_8x8bit m6036 (image[776],filter[6],mul_out[2012][25]);
mul_8x8bit m6037 (image[777],filter[7],mul_out[2012][26]);
mul_8x8bit m6038 (image[778],filter[8],mul_out[2012][27]);

adder_8bit ad670 (mul_out[2010][25],mul_out[2010][26],mul_out[2010][27],mul_out[2011][25],mul_out[2011][26],mul_out[2011][27],mul_out[2012][25],mul_out[2012][26],mul_out[2012][27],conv_out[670]);



mul_8x8bit m6039 (image[721],filter[0],mul_out[2013][25]);
mul_8x8bit m6040 (image[722],filter[1],mul_out[2013][26]);
mul_8x8bit m6041 (image[723],filter[2],mul_out[2013][27]);
mul_8x8bit m6042 (image[749],filter[3],mul_out[2014][25]);
mul_8x8bit m6043 (image[750],filter[4],mul_out[2014][26]);
mul_8x8bit m6044 (image[751],filter[5],mul_out[2014][27]);
mul_8x8bit m6045 (image[777],filter[6],mul_out[2015][25]);
mul_8x8bit m6046 (image[778],filter[7],mul_out[2015][26]);
mul_8x8bit m6047 (image[779],filter[8],mul_out[2015][27]);

adder_8bit ad671 (mul_out[2013][25],mul_out[2013][26],mul_out[2013][27],mul_out[2014][25],mul_out[2014][26],mul_out[2014][27],mul_out[2015][25],mul_out[2015][26],mul_out[2015][27],conv_out[671]);



mul_8x8bit m6048 (image[722],filter[0],mul_out[2016][25]);
mul_8x8bit m6049 (image[723],filter[1],mul_out[2016][26]);
mul_8x8bit m6050 (image[724],filter[2],mul_out[2016][27]);
mul_8x8bit m6051 (image[750],filter[3],mul_out[2017][25]);
mul_8x8bit m6052 (image[751],filter[4],mul_out[2017][26]);
mul_8x8bit m6053 (image[752],filter[5],mul_out[2017][27]);
mul_8x8bit m6054 (image[778],filter[6],mul_out[2018][25]);
mul_8x8bit m6055 (image[779],filter[7],mul_out[2018][26]);
mul_8x8bit m6056 (image[780],filter[8],mul_out[2018][27]);

adder_8bit ad672 (mul_out[2016][25],mul_out[2016][26],mul_out[2016][27],mul_out[2017][25],mul_out[2017][26],mul_out[2017][27],mul_out[2018][25],mul_out[2018][26],mul_out[2018][27],conv_out[672]);



mul_8x8bit m6057 (image[723],filter[0],mul_out[2019][25]);
mul_8x8bit m6058 (image[724],filter[1],mul_out[2019][26]);
mul_8x8bit m6059 (image[725],filter[2],mul_out[2019][27]);
mul_8x8bit m6060 (image[751],filter[3],mul_out[2020][25]);
mul_8x8bit m6061 (image[752],filter[4],mul_out[2020][26]);
mul_8x8bit m6062 (image[753],filter[5],mul_out[2020][27]);
mul_8x8bit m6063 (image[779],filter[6],mul_out[2021][25]);
mul_8x8bit m6064 (image[780],filter[7],mul_out[2021][26]);
mul_8x8bit m6065 (image[781],filter[8],mul_out[2021][27]);

adder_8bit ad673 (mul_out[2019][25],mul_out[2019][26],mul_out[2019][27],mul_out[2020][25],mul_out[2020][26],mul_out[2020][27],mul_out[2021][25],mul_out[2021][26],mul_out[2021][27],conv_out[673]);



mul_8x8bit m6066 (image[724],filter[0],mul_out[2022][25]);
mul_8x8bit m6067 (image[725],filter[1],mul_out[2022][26]);
mul_8x8bit m6068 (image[726],filter[2],mul_out[2022][27]);
mul_8x8bit m6069 (image[752],filter[3],mul_out[2023][25]);
mul_8x8bit m6070 (image[753],filter[4],mul_out[2023][26]);
mul_8x8bit m6071 (image[754],filter[5],mul_out[2023][27]);
mul_8x8bit m6072 (image[780],filter[6],mul_out[2024][25]);
mul_8x8bit m6073 (image[781],filter[7],mul_out[2024][26]);
mul_8x8bit m6074 (image[782],filter[8],mul_out[2024][27]);

adder_8bit ad674 (mul_out[2022][25],mul_out[2022][26],mul_out[2022][27],mul_out[2023][25],mul_out[2023][26],mul_out[2023][27],mul_out[2024][25],mul_out[2024][26],mul_out[2024][27],conv_out[674]);



mul_8x8bit m6075 (image[725],filter[0],mul_out[2025][25]);
mul_8x8bit m6076 (image[726],filter[1],mul_out[2025][26]);
mul_8x8bit m6077 (image[727],filter[2],mul_out[2025][27]);
mul_8x8bit m6078 (image[753],filter[3],mul_out[2026][25]);
mul_8x8bit m6079 (image[754],filter[4],mul_out[2026][26]);
mul_8x8bit m6080 (image[755],filter[5],mul_out[2026][27]);
mul_8x8bit m6081 (image[781],filter[6],mul_out[2027][25]);
mul_8x8bit m6082 (image[782],filter[7],mul_out[2027][26]);
mul_8x8bit m6083 (image[783],filter[8],mul_out[2027][27]);

adder_8bit ad675 (mul_out[2025][25],mul_out[2025][26],mul_out[2025][27],mul_out[2026][25],mul_out[2026][26],mul_out[2026][27],mul_out[2027][25],mul_out[2027][26],mul_out[2027][27],conv_out[675]);


endmodule



/* C code to generate above statements
// Online C compiler to run C program online
#include <stdio.h>

int main() {
   int d = 0;
 
   int k = 0;
   int l = 0;
   int n = 0;
    // Write C code here
    
int i = 0;




 int x = 0;
    for(int j = 0; j<26; j++){
      
      for(int i = 0; i<27; i++) {
        l = 0;
        if ((x+2) % 28 == 0) {
          x += 2;  
          continue;
      }     
      
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d,      x,      l,         k,   j);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+1,    x+1,      l+1,     k,   j+1);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+2,    x+2,      l+2,     k,   j+2);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+3,    x+28,    l+3,     k+1, j);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+4,    x+29,    l+4,   k+1, j+1);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+5,    x+30,    l+5,   k+1, j+2);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+6,    x+56,    l+6,     k+2, j);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n",d+7,    x+57,    l+7,   k+2, j+1);
    printf("mul_8x8bit m%d (image[%d],filter[%d],mul_out[%d][%d]);\n\n",d+8,  x+58,    l+8, k+2, j+2);
    
    printf("adder_8bit ad%d (mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],mul_out[%d][%d],conv_out[%d]);\n\n\n\n",n,k,j,k,j+1,k,j+2,k+1,j,k+1,j+1,k+1,j+2,k+2,j,k+2,j+1,k+2,j+2,n);
    
    n = n+1;
    k = k+3;
    
   //j = j+1;
    d =d +9;
    x = x+1;
  


   }
    }
   
    
    
    return 0;
}




*/
