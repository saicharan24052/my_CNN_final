`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/17/2025 02:31:40 PM
// Design Name: 
// Module Name: matrix_mul200x64
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module multi_7x28(// write the logic for MSB signed bit , includes the 2's COMPLIMENT module
input logic clk,rst,
input logic signed [8:0] mul_A,
input logic signed [32:0] mul_B,
output logic signed [40:0] mul_res

);

assign mul_res = mul_A*mul_B;

endmodule


module adder_200in (
input logic clk,rst,
 input logic signed [40:0] in_A_0,  
 input logic signed [40:0] in_A_1,   
 input logic signed [40:0] in_A_2,   
 input logic signed [40:0] in_A_3,   
 input logic signed [40:0] in_A_4,   
 input logic signed [40:0] in_A_5,   
 input logic signed [40:0] in_A_6,   
 input logic signed [40:0] in_A_7,   
 input logic signed [40:0] in_A_8,   
 input logic signed [40:0] in_A_9,   
 input logic signed [40:0] in_A_10,  
 input logic signed [40:0] in_A_11,  
 input logic signed [40:0] in_A_12,  
 input logic signed [40:0] in_A_13,  
 input logic signed [40:0] in_A_14,  
 input logic signed [40:0] in_A_15,  
 input logic signed [40:0] in_A_16,  
 input logic signed [40:0] in_A_17,  
 input logic signed [40:0] in_A_18,
 input logic signed [40:0] in_A_19,
 input logic signed [40:0] in_A_20,
 input logic signed [40:0] in_A_21,
 input logic signed [40:0] in_A_22,
 input logic signed [40:0] in_A_23,
 input logic signed [40:0] in_A_24,
 input logic signed [40:0] in_A_25,
 input logic signed [40:0] in_A_26,
 input logic signed [40:0] in_A_27,
 input logic signed [40:0] in_A_28,
 input logic signed [40:0] in_A_29,
 input logic signed [40:0] in_A_30,
 input logic signed [40:0] in_A_31,
 input logic signed [40:0] in_A_32,
 input logic signed [40:0] in_A_33,
 input logic signed [40:0] in_A_34,
 input logic signed [40:0] in_A_35,
 input logic signed [40:0] in_A_36,
 input logic signed [40:0] in_A_37,
 input logic signed [40:0] in_A_38,
 input logic signed [40:0] in_A_39,
 input logic signed [40:0] in_A_40,
 input logic signed [40:0] in_A_41,
 input logic signed [40:0] in_A_42,
 input logic signed [40:0] in_A_43,
 input logic signed [40:0] in_A_44,
 input logic signed [40:0] in_A_45,
 input logic signed [40:0] in_A_46,
 input logic signed [40:0] in_A_47,
 input logic signed [40:0] in_A_48,
 input logic signed [40:0] in_A_49,
 input logic signed [40:0] in_A_50,
 input logic signed [40:0] in_A_51,
 input logic signed [40:0] in_A_52,
 input logic signed [40:0] in_A_53,
 input logic signed [40:0] in_A_54,
 input logic signed [40:0] in_A_55,
 input logic signed [40:0] in_A_56,
 input logic signed [40:0] in_A_57,
 input logic signed [40:0] in_A_58,
 input logic signed [40:0] in_A_59,
 input logic signed [40:0] in_A_60,
 input logic signed [40:0] in_A_61,
 input logic signed [40:0] in_A_62,
 input logic signed [40:0] in_A_63,
 input logic signed [40:0] in_A_64,
 input logic signed [40:0] in_A_65,
 input logic signed [40:0] in_A_66,
 input logic signed [40:0] in_A_67,
 input logic signed [40:0] in_A_68,
 input logic signed [40:0] in_A_69,
 input logic signed [40:0] in_A_70,
 input logic signed [40:0] in_A_71,
 input logic signed [40:0] in_A_72,
 input logic signed [40:0] in_A_73,
 input logic signed [40:0] in_A_74,
 input logic signed [40:0] in_A_75,
 input logic signed [40:0] in_A_76,
 input logic signed [40:0] in_A_77,
 input logic signed [40:0] in_A_78,
 input logic signed [40:0] in_A_79,
 input logic signed [40:0] in_A_80,
 input logic signed [40:0] in_A_81,
 input logic signed [40:0] in_A_82,
 input logic signed [40:0] in_A_83,
 input logic signed [40:0] in_A_84,
 input logic signed [40:0] in_A_85,
 input logic signed [40:0] in_A_86,
 input logic signed [40:0] in_A_87,
 input logic signed [40:0] in_A_88,
 input logic signed [40:0] in_A_89,
 input logic signed [40:0] in_A_90,
 input logic signed [40:0] in_A_91,
 input logic signed [40:0] in_A_92,
 input logic signed [40:0] in_A_93,
 input logic signed [40:0] in_A_94,
 input logic signed [40:0] in_A_95,
 input logic signed [40:0] in_A_96,
 input logic signed [40:0] in_A_97,
 input logic signed [40:0] in_A_98,
 input logic signed [40:0] in_A_99,
 input logic signed [40:0] in_A_100,
 input logic signed [40:0] in_A_101,
 input logic signed [40:0] in_A_102,
 input logic signed [40:0] in_A_103,
 input logic signed [40:0] in_A_104,
 input logic signed [40:0] in_A_105,
 input logic signed [40:0] in_A_106,
 input logic signed [40:0] in_A_107,
 input logic signed [40:0] in_A_108,
 input logic signed [40:0] in_A_109,
 input logic signed [40:0] in_A_110,  
 input logic signed [40:0] in_A_111,
 input logic signed [40:0] in_A_112,
 input logic signed [40:0] in_A_113,
 input logic signed [40:0] in_A_114,
 input logic signed [40:0] in_A_115,
 input logic signed [40:0] in_A_116,
 input logic signed [40:0] in_A_117,
 input logic signed [40:0] in_A_118,
 input logic signed [40:0] in_A_119,
 input logic signed [40:0] in_A_120,
 input logic signed [40:0] in_A_121,
 input logic signed [40:0] in_A_122,
 input logic signed [40:0] in_A_123,
 input logic signed [40:0] in_A_124,
 input logic signed [40:0] in_A_125,
 input logic signed [40:0] in_A_126,
 input logic signed [40:0] in_A_127,
 input logic signed [40:0] in_A_128,
 input logic signed [40:0] in_A_129,
 input logic signed [40:0] in_A_130,
 input logic signed [40:0] in_A_131,
 input logic signed [40:0] in_A_132,
 input logic signed [40:0] in_A_133,
 input logic signed [40:0] in_A_134,
 input logic signed [40:0] in_A_135,
 input logic signed [40:0] in_A_136,
 input logic signed [40:0] in_A_137,
 input logic signed [40:0] in_A_138,
 input logic signed [40:0] in_A_139,
 input logic signed [40:0] in_A_140,
 input logic signed [40:0] in_A_141,
 input logic signed [40:0] in_A_142,
 input logic signed [40:0] in_A_143,
 input logic signed [40:0] in_A_144,
 input logic signed [40:0] in_A_145,
 input logic signed [40:0] in_A_146,
 input logic signed [40:0] in_A_147,
 input logic signed [40:0] in_A_148,
 input logic signed [40:0] in_A_149,
 input logic signed [40:0] in_A_150,
 input logic signed [40:0] in_A_151,
 input logic signed [40:0] in_A_152,
 input logic signed [40:0] in_A_153,
 input logic signed [40:0] in_A_154,
 input logic signed [40:0] in_A_155,
 input logic signed [40:0] in_A_156,
 input logic signed [40:0] in_A_157,
 input logic signed [40:0] in_A_158,
 input logic signed [40:0] in_A_159,
 input logic signed [40:0] in_A_160,
 input logic signed [40:0] in_A_161,
 input logic signed [40:0] in_A_162,
 input logic signed [40:0] in_A_163,
 input logic signed [40:0] in_A_164,
 input logic signed [40:0] in_A_165,
 input logic signed [40:0] in_A_166,
 input logic signed [40:0] in_A_167,
 input logic signed [40:0] in_A_168,
 input logic signed [40:0] in_A_169,
 input logic signed [40:0] in_A_170,
 input logic signed [40:0] in_A_171,
 input logic signed [40:0] in_A_172,
 input logic signed [40:0] in_A_173,
 input logic signed [40:0] in_A_174,
 input logic signed [40:0] in_A_175,
 input logic signed [40:0] in_A_176,
 input logic signed [40:0] in_A_177,
 input logic signed [40:0] in_A_178,
 input logic signed [40:0] in_A_179,
 input logic signed [40:0] in_A_180,
 input logic signed [40:0] in_A_181,
 input logic signed [40:0] in_A_182,
 input logic signed [40:0] in_A_183,
 input logic signed [40:0] in_A_184,
 input logic signed [40:0] in_A_185,
 input logic signed [40:0] in_A_186,
 input logic signed [40:0] in_A_187,
 input logic signed [40:0] in_A_188,
 input logic signed [40:0] in_A_189,
 input logic signed [40:0] in_A_190,
 input logic signed [40:0] in_A_191,
 input logic signed [40:0] in_A_192,
 input logic signed [40:0] in_A_193,
 input logic signed [40:0] in_A_194,
 input logic signed [40:0] in_A_195,
 input logic signed [40:0] in_A_196,
 input logic signed [40:0] in_A_197,
 input logic signed [40:0] in_A_198,
 input logic signed [40:0] in_A_199,
output logic signed  [47:0] out_A 
);

assign out_A = in_A_0 + in_A_1 + in_A_2 + in_A_3 + in_A_4 + in_A_5 + in_A_6 + in_A_7 + in_A_8 + in_A_9 + in_A_10 + in_A_11 + in_A_12 + in_A_13 + in_A_14 + in_A_15 + in_A_16 + in_A_17 + in_A_18 + in_A_19 + in_A_20 + in_A_21 + in_A_22 + in_A_23 + in_A_24 + in_A_25
 + in_A_26 + in_A_27 + in_A_28 + in_A_29 + in_A_30 + in_A_31 + in_A_32 + in_A_33 + in_A_34 + in_A_35 + in_A_36 + in_A_37 + in_A_38 + in_A_39 + in_A_40 + in_A_41 + in_A_42 + in_A_43 + in_A_44 + in_A_45 + in_A_46 + in_A_47 + in_A_48 + in_A_49 + in_A_50 + in_A_51 +
  in_A_52 + in_A_53 + in_A_54 + in_A_55 + in_A_56 + in_A_57 + in_A_58 + in_A_59 + in_A_60 + in_A_61 + in_A_62 + in_A_63 + in_A_64 + in_A_65 + in_A_66 + in_A_67 + in_A_68 + in_A_69 + in_A_70 + in_A_71 + in_A_72 + in_A_73 + in_A_74 + in_A_75 + in_A_76 + in_A_77 
+ in_A_78 + in_A_79 + in_A_80 + in_A_81 + in_A_82 + in_A_83 + in_A_84 + in_A_85 + in_A_86 + in_A_87 + in_A_88 + in_A_89 + in_A_90 + in_A_91 + in_A_92 + in_A_93 + in_A_94 + in_A_95 + in_A_96 + in_A_97 + in_A_98 + in_A_99 + in_A_100 + in_A_101 + in_A_102 + in_A_103
 + in_A_104 + in_A_105 + in_A_106 + in_A_107 + in_A_108 + in_A_109 + in_A_110 + in_A_111 + in_A_112 + in_A_113 + in_A_114 + in_A_115 + in_A_116 + in_A_117 + in_A_118 + in_A_119 + in_A_120 + in_A_121 + in_A_122 + in_A_123 + in_A_124 + in_A_125 + in_A_126 + in_A_127
  + in_A_128 + in_A_129 + in_A_130 + in_A_131 + in_A_132 + in_A_133 + in_A_134 + in_A_135 + in_A_136 + in_A_137 + in_A_138 + in_A_139 + in_A_140 + in_A_141 + in_A_142 + in_A_143 + in_A_144 + in_A_145 + in_A_146 + in_A_147 + in_A_148 + in_A_149 + in_A_150 + in_A_151
   + in_A_152 + in_A_153 + in_A_154 + in_A_155 + in_A_156 + in_A_157 + in_A_158 + in_A_159 + in_A_160 + in_A_161 + in_A_162 + in_A_163 + in_A_164 + in_A_165 + in_A_166 + in_A_167 + in_A_168 + in_A_169 + in_A_170 + in_A_171 + in_A_172 + in_A_173 + in_A_174 + in_A_175
    + in_A_176 + in_A_177 + in_A_178 + in_A_179 + in_A_180 + in_A_181 + in_A_182 + in_A_183 + in_A_184 + in_A_185 + in_A_186 + in_A_187 + in_A_188 + in_A_189 + in_A_190 + in_A_191 + in_A_192 + in_A_193 + in_A_194 + in_A_195 + in_A_196 + in_A_197 + in_A_198 + in_A_199;


endmodule



module matrix_mul200x64(  //actually 64 x 200
input logic clk,rst,
input logic signed [8:0]matrix_A [0:12799], //200*64
input logic signed [32:0]matrix_B [0:199], // flattened
output logic signed  [47:0] result_fc1[0:63]
    );
    
  
   
    
 logic signed [40:0] mul_res1 [0:12799];


multi_7x28 multi_7x28_mod_0(clk,rst,matrix_A[0],matrix_B[0],mul_res1[0]);
multi_7x28 multi_7x28_mod_1(clk,rst,matrix_A[1],matrix_B[1],mul_res1[1]);    
multi_7x28 multi_7x28_mod_2(clk,rst,matrix_A[2],matrix_B[2],mul_res1[2]);    
multi_7x28 multi_7x28_mod_3(clk,rst,matrix_A[3],matrix_B[3],mul_res1[3]);    
multi_7x28 multi_7x28_mod_4(clk,rst,matrix_A[4],matrix_B[4],mul_res1[4]);    
multi_7x28 multi_7x28_mod_5(clk,rst,matrix_A[5],matrix_B[5],mul_res1[5]);    
multi_7x28 multi_7x28_mod_6(clk,rst,matrix_A[6],matrix_B[6],mul_res1[6]);    
multi_7x28 multi_7x28_mod_7(clk,rst,matrix_A[7],matrix_B[7],mul_res1[7]);    
multi_7x28 multi_7x28_mod_8(clk,rst,matrix_A[8],matrix_B[8],mul_res1[8]);    
multi_7x28 multi_7x28_mod_9(clk,rst,matrix_A[9],matrix_B[9],mul_res1[9]);    
multi_7x28 multi_7x28_mod_10(clk,rst,matrix_A[10],matrix_B[10],mul_res1[10]);
multi_7x28 multi_7x28_mod_11(clk,rst,matrix_A[11],matrix_B[11],mul_res1[11]);
multi_7x28 multi_7x28_mod_12(clk,rst,matrix_A[12],matrix_B[12],mul_res1[12]);
multi_7x28 multi_7x28_mod_13(clk,rst,matrix_A[13],matrix_B[13],mul_res1[13]);
multi_7x28 multi_7x28_mod_14(clk,rst,matrix_A[14],matrix_B[14],mul_res1[14]);
multi_7x28 multi_7x28_mod_15(clk,rst,matrix_A[15],matrix_B[15],mul_res1[15]);
multi_7x28 multi_7x28_mod_16(clk,rst,matrix_A[16],matrix_B[16],mul_res1[16]);
multi_7x28 multi_7x28_mod_17(clk,rst,matrix_A[17],matrix_B[17],mul_res1[17]);
multi_7x28 multi_7x28_mod_18(clk,rst,matrix_A[18],matrix_B[18],mul_res1[18]);
multi_7x28 multi_7x28_mod_19(clk,rst,matrix_A[19],matrix_B[19],mul_res1[19]);
multi_7x28 multi_7x28_mod_20(clk,rst,matrix_A[20],matrix_B[20],mul_res1[20]);
multi_7x28 multi_7x28_mod_21(clk,rst,matrix_A[21],matrix_B[21],mul_res1[21]);
multi_7x28 multi_7x28_mod_22(clk,rst,matrix_A[22],matrix_B[22],mul_res1[22]);
multi_7x28 multi_7x28_mod_23(clk,rst,matrix_A[23],matrix_B[23],mul_res1[23]);
multi_7x28 multi_7x28_mod_24(clk,rst,matrix_A[24],matrix_B[24],mul_res1[24]);
multi_7x28 multi_7x28_mod_25(clk,rst,matrix_A[25],matrix_B[25],mul_res1[25]);
multi_7x28 multi_7x28_mod_26(clk,rst,matrix_A[26],matrix_B[26],mul_res1[26]);
multi_7x28 multi_7x28_mod_27(clk,rst,matrix_A[27],matrix_B[27],mul_res1[27]);
multi_7x28 multi_7x28_mod_28(clk,rst,matrix_A[28],matrix_B[28],mul_res1[28]);
multi_7x28 multi_7x28_mod_29(clk,rst,matrix_A[29],matrix_B[29],mul_res1[29]);
multi_7x28 multi_7x28_mod_30(clk,rst,matrix_A[30],matrix_B[30],mul_res1[30]);
multi_7x28 multi_7x28_mod_31(clk,rst,matrix_A[31],matrix_B[31],mul_res1[31]);
multi_7x28 multi_7x28_mod_32(clk,rst,matrix_A[32],matrix_B[32],mul_res1[32]);
multi_7x28 multi_7x28_mod_33(clk,rst,matrix_A[33],matrix_B[33],mul_res1[33]);
multi_7x28 multi_7x28_mod_34(clk,rst,matrix_A[34],matrix_B[34],mul_res1[34]);
multi_7x28 multi_7x28_mod_35(clk,rst,matrix_A[35],matrix_B[35],mul_res1[35]);
multi_7x28 multi_7x28_mod_36(clk,rst,matrix_A[36],matrix_B[36],mul_res1[36]);
multi_7x28 multi_7x28_mod_37(clk,rst,matrix_A[37],matrix_B[37],mul_res1[37]);
multi_7x28 multi_7x28_mod_38(clk,rst,matrix_A[38],matrix_B[38],mul_res1[38]);
multi_7x28 multi_7x28_mod_39(clk,rst,matrix_A[39],matrix_B[39],mul_res1[39]);
multi_7x28 multi_7x28_mod_40(clk,rst,matrix_A[40],matrix_B[40],mul_res1[40]);
multi_7x28 multi_7x28_mod_41(clk,rst,matrix_A[41],matrix_B[41],mul_res1[41]);
multi_7x28 multi_7x28_mod_42(clk,rst,matrix_A[42],matrix_B[42],mul_res1[42]);
multi_7x28 multi_7x28_mod_43(clk,rst,matrix_A[43],matrix_B[43],mul_res1[43]);
multi_7x28 multi_7x28_mod_44(clk,rst,matrix_A[44],matrix_B[44],mul_res1[44]);
multi_7x28 multi_7x28_mod_45(clk,rst,matrix_A[45],matrix_B[45],mul_res1[45]);
multi_7x28 multi_7x28_mod_46(clk,rst,matrix_A[46],matrix_B[46],mul_res1[46]);
multi_7x28 multi_7x28_mod_47(clk,rst,matrix_A[47],matrix_B[47],mul_res1[47]);
multi_7x28 multi_7x28_mod_48(clk,rst,matrix_A[48],matrix_B[48],mul_res1[48]);
multi_7x28 multi_7x28_mod_49(clk,rst,matrix_A[49],matrix_B[49],mul_res1[49]);
multi_7x28 multi_7x28_mod_50(clk,rst,matrix_A[50],matrix_B[50],mul_res1[50]);
multi_7x28 multi_7x28_mod_51(clk,rst,matrix_A[51],matrix_B[51],mul_res1[51]);
multi_7x28 multi_7x28_mod_52(clk,rst,matrix_A[52],matrix_B[52],mul_res1[52]);
multi_7x28 multi_7x28_mod_53(clk,rst,matrix_A[53],matrix_B[53],mul_res1[53]);
multi_7x28 multi_7x28_mod_54(clk,rst,matrix_A[54],matrix_B[54],mul_res1[54]);
multi_7x28 multi_7x28_mod_55(clk,rst,matrix_A[55],matrix_B[55],mul_res1[55]);
multi_7x28 multi_7x28_mod_56(clk,rst,matrix_A[56],matrix_B[56],mul_res1[56]);
multi_7x28 multi_7x28_mod_57(clk,rst,matrix_A[57],matrix_B[57],mul_res1[57]);
multi_7x28 multi_7x28_mod_58(clk,rst,matrix_A[58],matrix_B[58],mul_res1[58]);
multi_7x28 multi_7x28_mod_59(clk,rst,matrix_A[59],matrix_B[59],mul_res1[59]);
multi_7x28 multi_7x28_mod_60(clk,rst,matrix_A[60],matrix_B[60],mul_res1[60]);
multi_7x28 multi_7x28_mod_61(clk,rst,matrix_A[61],matrix_B[61],mul_res1[61]);
multi_7x28 multi_7x28_mod_62(clk,rst,matrix_A[62],matrix_B[62],mul_res1[62]);
multi_7x28 multi_7x28_mod_63(clk,rst,matrix_A[63],matrix_B[63],mul_res1[63]);
multi_7x28 multi_7x28_mod_64(clk,rst,matrix_A[64],matrix_B[64],mul_res1[64]);
multi_7x28 multi_7x28_mod_65(clk,rst,matrix_A[65],matrix_B[65],mul_res1[65]);
multi_7x28 multi_7x28_mod_66(clk,rst,matrix_A[66],matrix_B[66],mul_res1[66]);
multi_7x28 multi_7x28_mod_67(clk,rst,matrix_A[67],matrix_B[67],mul_res1[67]);
multi_7x28 multi_7x28_mod_68(clk,rst,matrix_A[68],matrix_B[68],mul_res1[68]);
multi_7x28 multi_7x28_mod_69(clk,rst,matrix_A[69],matrix_B[69],mul_res1[69]);
multi_7x28 multi_7x28_mod_70(clk,rst,matrix_A[70],matrix_B[70],mul_res1[70]);
multi_7x28 multi_7x28_mod_71(clk,rst,matrix_A[71],matrix_B[71],mul_res1[71]);
multi_7x28 multi_7x28_mod_72(clk,rst,matrix_A[72],matrix_B[72],mul_res1[72]);
multi_7x28 multi_7x28_mod_73(clk,rst,matrix_A[73],matrix_B[73],mul_res1[73]);
multi_7x28 multi_7x28_mod_74(clk,rst,matrix_A[74],matrix_B[74],mul_res1[74]);
multi_7x28 multi_7x28_mod_75(clk,rst,matrix_A[75],matrix_B[75],mul_res1[75]);
multi_7x28 multi_7x28_mod_76(clk,rst,matrix_A[76],matrix_B[76],mul_res1[76]);
multi_7x28 multi_7x28_mod_77(clk,rst,matrix_A[77],matrix_B[77],mul_res1[77]);
multi_7x28 multi_7x28_mod_78(clk,rst,matrix_A[78],matrix_B[78],mul_res1[78]);
multi_7x28 multi_7x28_mod_79(clk,rst,matrix_A[79],matrix_B[79],mul_res1[79]);
multi_7x28 multi_7x28_mod_80(clk,rst,matrix_A[80],matrix_B[80],mul_res1[80]);
multi_7x28 multi_7x28_mod_81(clk,rst,matrix_A[81],matrix_B[81],mul_res1[81]);
multi_7x28 multi_7x28_mod_82(clk,rst,matrix_A[82],matrix_B[82],mul_res1[82]);
multi_7x28 multi_7x28_mod_83(clk,rst,matrix_A[83],matrix_B[83],mul_res1[83]);
multi_7x28 multi_7x28_mod_84(clk,rst,matrix_A[84],matrix_B[84],mul_res1[84]);
multi_7x28 multi_7x28_mod_85(clk,rst,matrix_A[85],matrix_B[85],mul_res1[85]);
multi_7x28 multi_7x28_mod_86(clk,rst,matrix_A[86],matrix_B[86],mul_res1[86]);
multi_7x28 multi_7x28_mod_87(clk,rst,matrix_A[87],matrix_B[87],mul_res1[87]);
multi_7x28 multi_7x28_mod_88(clk,rst,matrix_A[88],matrix_B[88],mul_res1[88]);
multi_7x28 multi_7x28_mod_89(clk,rst,matrix_A[89],matrix_B[89],mul_res1[89]);
multi_7x28 multi_7x28_mod_90(clk,rst,matrix_A[90],matrix_B[90],mul_res1[90]);
multi_7x28 multi_7x28_mod_91(clk,rst,matrix_A[91],matrix_B[91],mul_res1[91]);
multi_7x28 multi_7x28_mod_92(clk,rst,matrix_A[92],matrix_B[92],mul_res1[92]);
multi_7x28 multi_7x28_mod_93(clk,rst,matrix_A[93],matrix_B[93],mul_res1[93]);
multi_7x28 multi_7x28_mod_94(clk,rst,matrix_A[94],matrix_B[94],mul_res1[94]);
multi_7x28 multi_7x28_mod_95(clk,rst,matrix_A[95],matrix_B[95],mul_res1[95]);
multi_7x28 multi_7x28_mod_96(clk,rst,matrix_A[96],matrix_B[96],mul_res1[96]);
multi_7x28 multi_7x28_mod_97(clk,rst,matrix_A[97],matrix_B[97],mul_res1[97]);
multi_7x28 multi_7x28_mod_98(clk,rst,matrix_A[98],matrix_B[98],mul_res1[98]);
multi_7x28 multi_7x28_mod_99(clk,rst,matrix_A[99],matrix_B[99],mul_res1[99]);
multi_7x28 multi_7x28_mod_100(clk,rst,matrix_A[100],matrix_B[100],mul_res1[100]);
multi_7x28 multi_7x28_mod_101(clk,rst,matrix_A[101],matrix_B[101],mul_res1[101]);
multi_7x28 multi_7x28_mod_102(clk,rst,matrix_A[102],matrix_B[102],mul_res1[102]);
multi_7x28 multi_7x28_mod_103(clk,rst,matrix_A[103],matrix_B[103],mul_res1[103]);
multi_7x28 multi_7x28_mod_104(clk,rst,matrix_A[104],matrix_B[104],mul_res1[104]);
multi_7x28 multi_7x28_mod_105(clk,rst,matrix_A[105],matrix_B[105],mul_res1[105]);
multi_7x28 multi_7x28_mod_106(clk,rst,matrix_A[106],matrix_B[106],mul_res1[106]);
multi_7x28 multi_7x28_mod_107(clk,rst,matrix_A[107],matrix_B[107],mul_res1[107]);
multi_7x28 multi_7x28_mod_108(clk,rst,matrix_A[108],matrix_B[108],mul_res1[108]);
multi_7x28 multi_7x28_mod_109(clk,rst,matrix_A[109],matrix_B[109],mul_res1[109]);
multi_7x28 multi_7x28_mod_110(clk,rst,matrix_A[110],matrix_B[110],mul_res1[110]);
multi_7x28 multi_7x28_mod_111(clk,rst,matrix_A[111],matrix_B[111],mul_res1[111]);
multi_7x28 multi_7x28_mod_112(clk,rst,matrix_A[112],matrix_B[112],mul_res1[112]);
multi_7x28 multi_7x28_mod_113(clk,rst,matrix_A[113],matrix_B[113],mul_res1[113]);
multi_7x28 multi_7x28_mod_114(clk,rst,matrix_A[114],matrix_B[114],mul_res1[114]);
multi_7x28 multi_7x28_mod_115(clk,rst,matrix_A[115],matrix_B[115],mul_res1[115]);
multi_7x28 multi_7x28_mod_116(clk,rst,matrix_A[116],matrix_B[116],mul_res1[116]);
multi_7x28 multi_7x28_mod_117(clk,rst,matrix_A[117],matrix_B[117],mul_res1[117]);
multi_7x28 multi_7x28_mod_118(clk,rst,matrix_A[118],matrix_B[118],mul_res1[118]);
multi_7x28 multi_7x28_mod_119(clk,rst,matrix_A[119],matrix_B[119],mul_res1[119]);
multi_7x28 multi_7x28_mod_120(clk,rst,matrix_A[120],matrix_B[120],mul_res1[120]);
multi_7x28 multi_7x28_mod_121(clk,rst,matrix_A[121],matrix_B[121],mul_res1[121]);
multi_7x28 multi_7x28_mod_122(clk,rst,matrix_A[122],matrix_B[122],mul_res1[122]);
multi_7x28 multi_7x28_mod_123(clk,rst,matrix_A[123],matrix_B[123],mul_res1[123]);
multi_7x28 multi_7x28_mod_124(clk,rst,matrix_A[124],matrix_B[124],mul_res1[124]);
multi_7x28 multi_7x28_mod_125(clk,rst,matrix_A[125],matrix_B[125],mul_res1[125]);
multi_7x28 multi_7x28_mod_126(clk,rst,matrix_A[126],matrix_B[126],mul_res1[126]);
multi_7x28 multi_7x28_mod_127(clk,rst,matrix_A[127],matrix_B[127],mul_res1[127]);
multi_7x28 multi_7x28_mod_128(clk,rst,matrix_A[128],matrix_B[128],mul_res1[128]);
multi_7x28 multi_7x28_mod_129(clk,rst,matrix_A[129],matrix_B[129],mul_res1[129]);
multi_7x28 multi_7x28_mod_130(clk,rst,matrix_A[130],matrix_B[130],mul_res1[130]);
multi_7x28 multi_7x28_mod_131(clk,rst,matrix_A[131],matrix_B[131],mul_res1[131]);
multi_7x28 multi_7x28_mod_132(clk,rst,matrix_A[132],matrix_B[132],mul_res1[132]);
multi_7x28 multi_7x28_mod_133(clk,rst,matrix_A[133],matrix_B[133],mul_res1[133]);
multi_7x28 multi_7x28_mod_134(clk,rst,matrix_A[134],matrix_B[134],mul_res1[134]);
multi_7x28 multi_7x28_mod_135(clk,rst,matrix_A[135],matrix_B[135],mul_res1[135]);
multi_7x28 multi_7x28_mod_136(clk,rst,matrix_A[136],matrix_B[136],mul_res1[136]);
multi_7x28 multi_7x28_mod_137(clk,rst,matrix_A[137],matrix_B[137],mul_res1[137]);
multi_7x28 multi_7x28_mod_138(clk,rst,matrix_A[138],matrix_B[138],mul_res1[138]);
multi_7x28 multi_7x28_mod_139(clk,rst,matrix_A[139],matrix_B[139],mul_res1[139]);
multi_7x28 multi_7x28_mod_140(clk,rst,matrix_A[140],matrix_B[140],mul_res1[140]);
multi_7x28 multi_7x28_mod_141(clk,rst,matrix_A[141],matrix_B[141],mul_res1[141]);
multi_7x28 multi_7x28_mod_142(clk,rst,matrix_A[142],matrix_B[142],mul_res1[142]);
multi_7x28 multi_7x28_mod_143(clk,rst,matrix_A[143],matrix_B[143],mul_res1[143]);
multi_7x28 multi_7x28_mod_144(clk,rst,matrix_A[144],matrix_B[144],mul_res1[144]);
multi_7x28 multi_7x28_mod_145(clk,rst,matrix_A[145],matrix_B[145],mul_res1[145]);
multi_7x28 multi_7x28_mod_146(clk,rst,matrix_A[146],matrix_B[146],mul_res1[146]);
multi_7x28 multi_7x28_mod_147(clk,rst,matrix_A[147],matrix_B[147],mul_res1[147]);
multi_7x28 multi_7x28_mod_148(clk,rst,matrix_A[148],matrix_B[148],mul_res1[148]);
multi_7x28 multi_7x28_mod_149(clk,rst,matrix_A[149],matrix_B[149],mul_res1[149]);
multi_7x28 multi_7x28_mod_150(clk,rst,matrix_A[150],matrix_B[150],mul_res1[150]);
multi_7x28 multi_7x28_mod_151(clk,rst,matrix_A[151],matrix_B[151],mul_res1[151]);
multi_7x28 multi_7x28_mod_152(clk,rst,matrix_A[152],matrix_B[152],mul_res1[152]);
multi_7x28 multi_7x28_mod_153(clk,rst,matrix_A[153],matrix_B[153],mul_res1[153]);
multi_7x28 multi_7x28_mod_154(clk,rst,matrix_A[154],matrix_B[154],mul_res1[154]);
multi_7x28 multi_7x28_mod_155(clk,rst,matrix_A[155],matrix_B[155],mul_res1[155]);
multi_7x28 multi_7x28_mod_156(clk,rst,matrix_A[156],matrix_B[156],mul_res1[156]);
multi_7x28 multi_7x28_mod_157(clk,rst,matrix_A[157],matrix_B[157],mul_res1[157]);
multi_7x28 multi_7x28_mod_158(clk,rst,matrix_A[158],matrix_B[158],mul_res1[158]);
multi_7x28 multi_7x28_mod_159(clk,rst,matrix_A[159],matrix_B[159],mul_res1[159]);
multi_7x28 multi_7x28_mod_160(clk,rst,matrix_A[160],matrix_B[160],mul_res1[160]);
multi_7x28 multi_7x28_mod_161(clk,rst,matrix_A[161],matrix_B[161],mul_res1[161]);
multi_7x28 multi_7x28_mod_162(clk,rst,matrix_A[162],matrix_B[162],mul_res1[162]);
multi_7x28 multi_7x28_mod_163(clk,rst,matrix_A[163],matrix_B[163],mul_res1[163]);
multi_7x28 multi_7x28_mod_164(clk,rst,matrix_A[164],matrix_B[164],mul_res1[164]);
multi_7x28 multi_7x28_mod_165(clk,rst,matrix_A[165],matrix_B[165],mul_res1[165]);
multi_7x28 multi_7x28_mod_166(clk,rst,matrix_A[166],matrix_B[166],mul_res1[166]);
multi_7x28 multi_7x28_mod_167(clk,rst,matrix_A[167],matrix_B[167],mul_res1[167]);
multi_7x28 multi_7x28_mod_168(clk,rst,matrix_A[168],matrix_B[168],mul_res1[168]);
multi_7x28 multi_7x28_mod_169(clk,rst,matrix_A[169],matrix_B[169],mul_res1[169]);
multi_7x28 multi_7x28_mod_170(clk,rst,matrix_A[170],matrix_B[170],mul_res1[170]);
multi_7x28 multi_7x28_mod_171(clk,rst,matrix_A[171],matrix_B[171],mul_res1[171]);
multi_7x28 multi_7x28_mod_172(clk,rst,matrix_A[172],matrix_B[172],mul_res1[172]);
multi_7x28 multi_7x28_mod_173(clk,rst,matrix_A[173],matrix_B[173],mul_res1[173]);
multi_7x28 multi_7x28_mod_174(clk,rst,matrix_A[174],matrix_B[174],mul_res1[174]);
multi_7x28 multi_7x28_mod_175(clk,rst,matrix_A[175],matrix_B[175],mul_res1[175]);
multi_7x28 multi_7x28_mod_176(clk,rst,matrix_A[176],matrix_B[176],mul_res1[176]);
multi_7x28 multi_7x28_mod_177(clk,rst,matrix_A[177],matrix_B[177],mul_res1[177]);
multi_7x28 multi_7x28_mod_178(clk,rst,matrix_A[178],matrix_B[178],mul_res1[178]);
multi_7x28 multi_7x28_mod_179(clk,rst,matrix_A[179],matrix_B[179],mul_res1[179]);
multi_7x28 multi_7x28_mod_180(clk,rst,matrix_A[180],matrix_B[180],mul_res1[180]);
multi_7x28 multi_7x28_mod_181(clk,rst,matrix_A[181],matrix_B[181],mul_res1[181]);
multi_7x28 multi_7x28_mod_182(clk,rst,matrix_A[182],matrix_B[182],mul_res1[182]);
multi_7x28 multi_7x28_mod_183(clk,rst,matrix_A[183],matrix_B[183],mul_res1[183]);
multi_7x28 multi_7x28_mod_184(clk,rst,matrix_A[184],matrix_B[184],mul_res1[184]);
multi_7x28 multi_7x28_mod_185(clk,rst,matrix_A[185],matrix_B[185],mul_res1[185]);
multi_7x28 multi_7x28_mod_186(clk,rst,matrix_A[186],matrix_B[186],mul_res1[186]);
multi_7x28 multi_7x28_mod_187(clk,rst,matrix_A[187],matrix_B[187],mul_res1[187]);
multi_7x28 multi_7x28_mod_188(clk,rst,matrix_A[188],matrix_B[188],mul_res1[188]);
multi_7x28 multi_7x28_mod_189(clk,rst,matrix_A[189],matrix_B[189],mul_res1[189]);
multi_7x28 multi_7x28_mod_190(clk,rst,matrix_A[190],matrix_B[190],mul_res1[190]);
multi_7x28 multi_7x28_mod_191(clk,rst,matrix_A[191],matrix_B[191],mul_res1[191]);
multi_7x28 multi_7x28_mod_192(clk,rst,matrix_A[192],matrix_B[192],mul_res1[192]);
multi_7x28 multi_7x28_mod_193(clk,rst,matrix_A[193],matrix_B[193],mul_res1[193]);
multi_7x28 multi_7x28_mod_194(clk,rst,matrix_A[194],matrix_B[194],mul_res1[194]);
multi_7x28 multi_7x28_mod_195(clk,rst,matrix_A[195],matrix_B[195],mul_res1[195]);
multi_7x28 multi_7x28_mod_196(clk,rst,matrix_A[196],matrix_B[196],mul_res1[196]);
multi_7x28 multi_7x28_mod_197(clk,rst,matrix_A[197],matrix_B[197],mul_res1[197]);
multi_7x28 multi_7x28_mod_198(clk,rst,matrix_A[198],matrix_B[198],mul_res1[198]);
multi_7x28 multi_7x28_mod_199(clk,rst,matrix_A[199],matrix_B[199],mul_res1[199]);
multi_7x28 multi_7x28_mod_200(clk,rst,matrix_A[200],matrix_B[0],mul_res1[200]);
multi_7x28 multi_7x28_mod_201(clk,rst,matrix_A[201],matrix_B[1],mul_res1[201]);
multi_7x28 multi_7x28_mod_202(clk,rst,matrix_A[202],matrix_B[2],mul_res1[202]);
multi_7x28 multi_7x28_mod_203(clk,rst,matrix_A[203],matrix_B[3],mul_res1[203]);
multi_7x28 multi_7x28_mod_204(clk,rst,matrix_A[204],matrix_B[4],mul_res1[204]);
multi_7x28 multi_7x28_mod_205(clk,rst,matrix_A[205],matrix_B[5],mul_res1[205]);
multi_7x28 multi_7x28_mod_206(clk,rst,matrix_A[206],matrix_B[6],mul_res1[206]);
multi_7x28 multi_7x28_mod_207(clk,rst,matrix_A[207],matrix_B[7],mul_res1[207]);
multi_7x28 multi_7x28_mod_208(clk,rst,matrix_A[208],matrix_B[8],mul_res1[208]);
multi_7x28 multi_7x28_mod_209(clk,rst,matrix_A[209],matrix_B[9],mul_res1[209]);
multi_7x28 multi_7x28_mod_210(clk,rst,matrix_A[210],matrix_B[10],mul_res1[210]);
multi_7x28 multi_7x28_mod_211(clk,rst,matrix_A[211],matrix_B[11],mul_res1[211]);
multi_7x28 multi_7x28_mod_212(clk,rst,matrix_A[212],matrix_B[12],mul_res1[212]);
multi_7x28 multi_7x28_mod_213(clk,rst,matrix_A[213],matrix_B[13],mul_res1[213]);
multi_7x28 multi_7x28_mod_214(clk,rst,matrix_A[214],matrix_B[14],mul_res1[214]);
multi_7x28 multi_7x28_mod_215(clk,rst,matrix_A[215],matrix_B[15],mul_res1[215]);
multi_7x28 multi_7x28_mod_216(clk,rst,matrix_A[216],matrix_B[16],mul_res1[216]);
multi_7x28 multi_7x28_mod_217(clk,rst,matrix_A[217],matrix_B[17],mul_res1[217]);
multi_7x28 multi_7x28_mod_218(clk,rst,matrix_A[218],matrix_B[18],mul_res1[218]);
multi_7x28 multi_7x28_mod_219(clk,rst,matrix_A[219],matrix_B[19],mul_res1[219]);
multi_7x28 multi_7x28_mod_220(clk,rst,matrix_A[220],matrix_B[20],mul_res1[220]);
multi_7x28 multi_7x28_mod_221(clk,rst,matrix_A[221],matrix_B[21],mul_res1[221]);
multi_7x28 multi_7x28_mod_222(clk,rst,matrix_A[222],matrix_B[22],mul_res1[222]);
multi_7x28 multi_7x28_mod_223(clk,rst,matrix_A[223],matrix_B[23],mul_res1[223]);
multi_7x28 multi_7x28_mod_224(clk,rst,matrix_A[224],matrix_B[24],mul_res1[224]);
multi_7x28 multi_7x28_mod_225(clk,rst,matrix_A[225],matrix_B[25],mul_res1[225]);
multi_7x28 multi_7x28_mod_226(clk,rst,matrix_A[226],matrix_B[26],mul_res1[226]);
multi_7x28 multi_7x28_mod_227(clk,rst,matrix_A[227],matrix_B[27],mul_res1[227]);
multi_7x28 multi_7x28_mod_228(clk,rst,matrix_A[228],matrix_B[28],mul_res1[228]);
multi_7x28 multi_7x28_mod_229(clk,rst,matrix_A[229],matrix_B[29],mul_res1[229]);
multi_7x28 multi_7x28_mod_230(clk,rst,matrix_A[230],matrix_B[30],mul_res1[230]);
multi_7x28 multi_7x28_mod_231(clk,rst,matrix_A[231],matrix_B[31],mul_res1[231]);
multi_7x28 multi_7x28_mod_232(clk,rst,matrix_A[232],matrix_B[32],mul_res1[232]);
multi_7x28 multi_7x28_mod_233(clk,rst,matrix_A[233],matrix_B[33],mul_res1[233]);
multi_7x28 multi_7x28_mod_234(clk,rst,matrix_A[234],matrix_B[34],mul_res1[234]);
multi_7x28 multi_7x28_mod_235(clk,rst,matrix_A[235],matrix_B[35],mul_res1[235]);
multi_7x28 multi_7x28_mod_236(clk,rst,matrix_A[236],matrix_B[36],mul_res1[236]);
multi_7x28 multi_7x28_mod_237(clk,rst,matrix_A[237],matrix_B[37],mul_res1[237]);
multi_7x28 multi_7x28_mod_238(clk,rst,matrix_A[238],matrix_B[38],mul_res1[238]);
multi_7x28 multi_7x28_mod_239(clk,rst,matrix_A[239],matrix_B[39],mul_res1[239]);
multi_7x28 multi_7x28_mod_240(clk,rst,matrix_A[240],matrix_B[40],mul_res1[240]);
multi_7x28 multi_7x28_mod_241(clk,rst,matrix_A[241],matrix_B[41],mul_res1[241]);
multi_7x28 multi_7x28_mod_242(clk,rst,matrix_A[242],matrix_B[42],mul_res1[242]);
multi_7x28 multi_7x28_mod_243(clk,rst,matrix_A[243],matrix_B[43],mul_res1[243]);
multi_7x28 multi_7x28_mod_244(clk,rst,matrix_A[244],matrix_B[44],mul_res1[244]);
multi_7x28 multi_7x28_mod_245(clk,rst,matrix_A[245],matrix_B[45],mul_res1[245]);
multi_7x28 multi_7x28_mod_246(clk,rst,matrix_A[246],matrix_B[46],mul_res1[246]);
multi_7x28 multi_7x28_mod_247(clk,rst,matrix_A[247],matrix_B[47],mul_res1[247]);
multi_7x28 multi_7x28_mod_248(clk,rst,matrix_A[248],matrix_B[48],mul_res1[248]);
multi_7x28 multi_7x28_mod_249(clk,rst,matrix_A[249],matrix_B[49],mul_res1[249]);
multi_7x28 multi_7x28_mod_250(clk,rst,matrix_A[250],matrix_B[50],mul_res1[250]);
multi_7x28 multi_7x28_mod_251(clk,rst,matrix_A[251],matrix_B[51],mul_res1[251]);
multi_7x28 multi_7x28_mod_252(clk,rst,matrix_A[252],matrix_B[52],mul_res1[252]);
multi_7x28 multi_7x28_mod_253(clk,rst,matrix_A[253],matrix_B[53],mul_res1[253]);
multi_7x28 multi_7x28_mod_254(clk,rst,matrix_A[254],matrix_B[54],mul_res1[254]);
multi_7x28 multi_7x28_mod_255(clk,rst,matrix_A[255],matrix_B[55],mul_res1[255]);
multi_7x28 multi_7x28_mod_256(clk,rst,matrix_A[256],matrix_B[56],mul_res1[256]);
multi_7x28 multi_7x28_mod_257(clk,rst,matrix_A[257],matrix_B[57],mul_res1[257]);
multi_7x28 multi_7x28_mod_258(clk,rst,matrix_A[258],matrix_B[58],mul_res1[258]);
multi_7x28 multi_7x28_mod_259(clk,rst,matrix_A[259],matrix_B[59],mul_res1[259]);
multi_7x28 multi_7x28_mod_260(clk,rst,matrix_A[260],matrix_B[60],mul_res1[260]);
multi_7x28 multi_7x28_mod_261(clk,rst,matrix_A[261],matrix_B[61],mul_res1[261]);
multi_7x28 multi_7x28_mod_262(clk,rst,matrix_A[262],matrix_B[62],mul_res1[262]);
multi_7x28 multi_7x28_mod_263(clk,rst,matrix_A[263],matrix_B[63],mul_res1[263]);
multi_7x28 multi_7x28_mod_264(clk,rst,matrix_A[264],matrix_B[64],mul_res1[264]);
multi_7x28 multi_7x28_mod_265(clk,rst,matrix_A[265],matrix_B[65],mul_res1[265]);
multi_7x28 multi_7x28_mod_266(clk,rst,matrix_A[266],matrix_B[66],mul_res1[266]);
multi_7x28 multi_7x28_mod_267(clk,rst,matrix_A[267],matrix_B[67],mul_res1[267]);
multi_7x28 multi_7x28_mod_268(clk,rst,matrix_A[268],matrix_B[68],mul_res1[268]);
multi_7x28 multi_7x28_mod_269(clk,rst,matrix_A[269],matrix_B[69],mul_res1[269]);
multi_7x28 multi_7x28_mod_270(clk,rst,matrix_A[270],matrix_B[70],mul_res1[270]);
multi_7x28 multi_7x28_mod_271(clk,rst,matrix_A[271],matrix_B[71],mul_res1[271]);
multi_7x28 multi_7x28_mod_272(clk,rst,matrix_A[272],matrix_B[72],mul_res1[272]);
multi_7x28 multi_7x28_mod_273(clk,rst,matrix_A[273],matrix_B[73],mul_res1[273]);
multi_7x28 multi_7x28_mod_274(clk,rst,matrix_A[274],matrix_B[74],mul_res1[274]);
multi_7x28 multi_7x28_mod_275(clk,rst,matrix_A[275],matrix_B[75],mul_res1[275]);
multi_7x28 multi_7x28_mod_276(clk,rst,matrix_A[276],matrix_B[76],mul_res1[276]);
multi_7x28 multi_7x28_mod_277(clk,rst,matrix_A[277],matrix_B[77],mul_res1[277]);
multi_7x28 multi_7x28_mod_278(clk,rst,matrix_A[278],matrix_B[78],mul_res1[278]);
multi_7x28 multi_7x28_mod_279(clk,rst,matrix_A[279],matrix_B[79],mul_res1[279]);
multi_7x28 multi_7x28_mod_280(clk,rst,matrix_A[280],matrix_B[80],mul_res1[280]);
multi_7x28 multi_7x28_mod_281(clk,rst,matrix_A[281],matrix_B[81],mul_res1[281]);
multi_7x28 multi_7x28_mod_282(clk,rst,matrix_A[282],matrix_B[82],mul_res1[282]);
multi_7x28 multi_7x28_mod_283(clk,rst,matrix_A[283],matrix_B[83],mul_res1[283]);
multi_7x28 multi_7x28_mod_284(clk,rst,matrix_A[284],matrix_B[84],mul_res1[284]);
multi_7x28 multi_7x28_mod_285(clk,rst,matrix_A[285],matrix_B[85],mul_res1[285]);
multi_7x28 multi_7x28_mod_286(clk,rst,matrix_A[286],matrix_B[86],mul_res1[286]);
multi_7x28 multi_7x28_mod_287(clk,rst,matrix_A[287],matrix_B[87],mul_res1[287]);
multi_7x28 multi_7x28_mod_288(clk,rst,matrix_A[288],matrix_B[88],mul_res1[288]);
multi_7x28 multi_7x28_mod_289(clk,rst,matrix_A[289],matrix_B[89],mul_res1[289]);
multi_7x28 multi_7x28_mod_290(clk,rst,matrix_A[290],matrix_B[90],mul_res1[290]);
multi_7x28 multi_7x28_mod_291(clk,rst,matrix_A[291],matrix_B[91],mul_res1[291]);
multi_7x28 multi_7x28_mod_292(clk,rst,matrix_A[292],matrix_B[92],mul_res1[292]);
multi_7x28 multi_7x28_mod_293(clk,rst,matrix_A[293],matrix_B[93],mul_res1[293]);
multi_7x28 multi_7x28_mod_294(clk,rst,matrix_A[294],matrix_B[94],mul_res1[294]);
multi_7x28 multi_7x28_mod_295(clk,rst,matrix_A[295],matrix_B[95],mul_res1[295]);
multi_7x28 multi_7x28_mod_296(clk,rst,matrix_A[296],matrix_B[96],mul_res1[296]);
multi_7x28 multi_7x28_mod_297(clk,rst,matrix_A[297],matrix_B[97],mul_res1[297]);
multi_7x28 multi_7x28_mod_298(clk,rst,matrix_A[298],matrix_B[98],mul_res1[298]);
multi_7x28 multi_7x28_mod_299(clk,rst,matrix_A[299],matrix_B[99],mul_res1[299]);
multi_7x28 multi_7x28_mod_300(clk,rst,matrix_A[300],matrix_B[100],mul_res1[300]);
multi_7x28 multi_7x28_mod_301(clk,rst,matrix_A[301],matrix_B[101],mul_res1[301]);
multi_7x28 multi_7x28_mod_302(clk,rst,matrix_A[302],matrix_B[102],mul_res1[302]);
multi_7x28 multi_7x28_mod_303(clk,rst,matrix_A[303],matrix_B[103],mul_res1[303]);
multi_7x28 multi_7x28_mod_304(clk,rst,matrix_A[304],matrix_B[104],mul_res1[304]);
multi_7x28 multi_7x28_mod_305(clk,rst,matrix_A[305],matrix_B[105],mul_res1[305]);
multi_7x28 multi_7x28_mod_306(clk,rst,matrix_A[306],matrix_B[106],mul_res1[306]);
multi_7x28 multi_7x28_mod_307(clk,rst,matrix_A[307],matrix_B[107],mul_res1[307]);
multi_7x28 multi_7x28_mod_308(clk,rst,matrix_A[308],matrix_B[108],mul_res1[308]);
multi_7x28 multi_7x28_mod_309(clk,rst,matrix_A[309],matrix_B[109],mul_res1[309]);
multi_7x28 multi_7x28_mod_310(clk,rst,matrix_A[310],matrix_B[110],mul_res1[310]);
multi_7x28 multi_7x28_mod_311(clk,rst,matrix_A[311],matrix_B[111],mul_res1[311]);
multi_7x28 multi_7x28_mod_312(clk,rst,matrix_A[312],matrix_B[112],mul_res1[312]);
multi_7x28 multi_7x28_mod_313(clk,rst,matrix_A[313],matrix_B[113],mul_res1[313]);
multi_7x28 multi_7x28_mod_314(clk,rst,matrix_A[314],matrix_B[114],mul_res1[314]);
multi_7x28 multi_7x28_mod_315(clk,rst,matrix_A[315],matrix_B[115],mul_res1[315]);
multi_7x28 multi_7x28_mod_316(clk,rst,matrix_A[316],matrix_B[116],mul_res1[316]);
multi_7x28 multi_7x28_mod_317(clk,rst,matrix_A[317],matrix_B[117],mul_res1[317]);
multi_7x28 multi_7x28_mod_318(clk,rst,matrix_A[318],matrix_B[118],mul_res1[318]);
multi_7x28 multi_7x28_mod_319(clk,rst,matrix_A[319],matrix_B[119],mul_res1[319]);
multi_7x28 multi_7x28_mod_320(clk,rst,matrix_A[320],matrix_B[120],mul_res1[320]);
multi_7x28 multi_7x28_mod_321(clk,rst,matrix_A[321],matrix_B[121],mul_res1[321]);
multi_7x28 multi_7x28_mod_322(clk,rst,matrix_A[322],matrix_B[122],mul_res1[322]);
multi_7x28 multi_7x28_mod_323(clk,rst,matrix_A[323],matrix_B[123],mul_res1[323]);
multi_7x28 multi_7x28_mod_324(clk,rst,matrix_A[324],matrix_B[124],mul_res1[324]);
multi_7x28 multi_7x28_mod_325(clk,rst,matrix_A[325],matrix_B[125],mul_res1[325]);
multi_7x28 multi_7x28_mod_326(clk,rst,matrix_A[326],matrix_B[126],mul_res1[326]);
multi_7x28 multi_7x28_mod_327(clk,rst,matrix_A[327],matrix_B[127],mul_res1[327]);
multi_7x28 multi_7x28_mod_328(clk,rst,matrix_A[328],matrix_B[128],mul_res1[328]);
multi_7x28 multi_7x28_mod_329(clk,rst,matrix_A[329],matrix_B[129],mul_res1[329]);
multi_7x28 multi_7x28_mod_330(clk,rst,matrix_A[330],matrix_B[130],mul_res1[330]);
multi_7x28 multi_7x28_mod_331(clk,rst,matrix_A[331],matrix_B[131],mul_res1[331]);
multi_7x28 multi_7x28_mod_332(clk,rst,matrix_A[332],matrix_B[132],mul_res1[332]);
multi_7x28 multi_7x28_mod_333(clk,rst,matrix_A[333],matrix_B[133],mul_res1[333]);
multi_7x28 multi_7x28_mod_334(clk,rst,matrix_A[334],matrix_B[134],mul_res1[334]);
multi_7x28 multi_7x28_mod_335(clk,rst,matrix_A[335],matrix_B[135],mul_res1[335]);
multi_7x28 multi_7x28_mod_336(clk,rst,matrix_A[336],matrix_B[136],mul_res1[336]);
multi_7x28 multi_7x28_mod_337(clk,rst,matrix_A[337],matrix_B[137],mul_res1[337]);
multi_7x28 multi_7x28_mod_338(clk,rst,matrix_A[338],matrix_B[138],mul_res1[338]);
multi_7x28 multi_7x28_mod_339(clk,rst,matrix_A[339],matrix_B[139],mul_res1[339]);
multi_7x28 multi_7x28_mod_340(clk,rst,matrix_A[340],matrix_B[140],mul_res1[340]);
multi_7x28 multi_7x28_mod_341(clk,rst,matrix_A[341],matrix_B[141],mul_res1[341]);
multi_7x28 multi_7x28_mod_342(clk,rst,matrix_A[342],matrix_B[142],mul_res1[342]);
multi_7x28 multi_7x28_mod_343(clk,rst,matrix_A[343],matrix_B[143],mul_res1[343]);
multi_7x28 multi_7x28_mod_344(clk,rst,matrix_A[344],matrix_B[144],mul_res1[344]);
multi_7x28 multi_7x28_mod_345(clk,rst,matrix_A[345],matrix_B[145],mul_res1[345]);
multi_7x28 multi_7x28_mod_346(clk,rst,matrix_A[346],matrix_B[146],mul_res1[346]);
multi_7x28 multi_7x28_mod_347(clk,rst,matrix_A[347],matrix_B[147],mul_res1[347]);
multi_7x28 multi_7x28_mod_348(clk,rst,matrix_A[348],matrix_B[148],mul_res1[348]);
multi_7x28 multi_7x28_mod_349(clk,rst,matrix_A[349],matrix_B[149],mul_res1[349]);
multi_7x28 multi_7x28_mod_350(clk,rst,matrix_A[350],matrix_B[150],mul_res1[350]);
multi_7x28 multi_7x28_mod_351(clk,rst,matrix_A[351],matrix_B[151],mul_res1[351]);
multi_7x28 multi_7x28_mod_352(clk,rst,matrix_A[352],matrix_B[152],mul_res1[352]);
multi_7x28 multi_7x28_mod_353(clk,rst,matrix_A[353],matrix_B[153],mul_res1[353]);
multi_7x28 multi_7x28_mod_354(clk,rst,matrix_A[354],matrix_B[154],mul_res1[354]);
multi_7x28 multi_7x28_mod_355(clk,rst,matrix_A[355],matrix_B[155],mul_res1[355]);
multi_7x28 multi_7x28_mod_356(clk,rst,matrix_A[356],matrix_B[156],mul_res1[356]);
multi_7x28 multi_7x28_mod_357(clk,rst,matrix_A[357],matrix_B[157],mul_res1[357]);
multi_7x28 multi_7x28_mod_358(clk,rst,matrix_A[358],matrix_B[158],mul_res1[358]);
multi_7x28 multi_7x28_mod_359(clk,rst,matrix_A[359],matrix_B[159],mul_res1[359]);
multi_7x28 multi_7x28_mod_360(clk,rst,matrix_A[360],matrix_B[160],mul_res1[360]);
multi_7x28 multi_7x28_mod_361(clk,rst,matrix_A[361],matrix_B[161],mul_res1[361]);
multi_7x28 multi_7x28_mod_362(clk,rst,matrix_A[362],matrix_B[162],mul_res1[362]);
multi_7x28 multi_7x28_mod_363(clk,rst,matrix_A[363],matrix_B[163],mul_res1[363]);
multi_7x28 multi_7x28_mod_364(clk,rst,matrix_A[364],matrix_B[164],mul_res1[364]);
multi_7x28 multi_7x28_mod_365(clk,rst,matrix_A[365],matrix_B[165],mul_res1[365]);
multi_7x28 multi_7x28_mod_366(clk,rst,matrix_A[366],matrix_B[166],mul_res1[366]);
multi_7x28 multi_7x28_mod_367(clk,rst,matrix_A[367],matrix_B[167],mul_res1[367]);
multi_7x28 multi_7x28_mod_368(clk,rst,matrix_A[368],matrix_B[168],mul_res1[368]);
multi_7x28 multi_7x28_mod_369(clk,rst,matrix_A[369],matrix_B[169],mul_res1[369]);
multi_7x28 multi_7x28_mod_370(clk,rst,matrix_A[370],matrix_B[170],mul_res1[370]);
multi_7x28 multi_7x28_mod_371(clk,rst,matrix_A[371],matrix_B[171],mul_res1[371]);
multi_7x28 multi_7x28_mod_372(clk,rst,matrix_A[372],matrix_B[172],mul_res1[372]);
multi_7x28 multi_7x28_mod_373(clk,rst,matrix_A[373],matrix_B[173],mul_res1[373]);
multi_7x28 multi_7x28_mod_374(clk,rst,matrix_A[374],matrix_B[174],mul_res1[374]);
multi_7x28 multi_7x28_mod_375(clk,rst,matrix_A[375],matrix_B[175],mul_res1[375]);
multi_7x28 multi_7x28_mod_376(clk,rst,matrix_A[376],matrix_B[176],mul_res1[376]);
multi_7x28 multi_7x28_mod_377(clk,rst,matrix_A[377],matrix_B[177],mul_res1[377]);
multi_7x28 multi_7x28_mod_378(clk,rst,matrix_A[378],matrix_B[178],mul_res1[378]);
multi_7x28 multi_7x28_mod_379(clk,rst,matrix_A[379],matrix_B[179],mul_res1[379]);
multi_7x28 multi_7x28_mod_380(clk,rst,matrix_A[380],matrix_B[180],mul_res1[380]);
multi_7x28 multi_7x28_mod_381(clk,rst,matrix_A[381],matrix_B[181],mul_res1[381]);
multi_7x28 multi_7x28_mod_382(clk,rst,matrix_A[382],matrix_B[182],mul_res1[382]);
multi_7x28 multi_7x28_mod_383(clk,rst,matrix_A[383],matrix_B[183],mul_res1[383]);
multi_7x28 multi_7x28_mod_384(clk,rst,matrix_A[384],matrix_B[184],mul_res1[384]);
multi_7x28 multi_7x28_mod_385(clk,rst,matrix_A[385],matrix_B[185],mul_res1[385]);
multi_7x28 multi_7x28_mod_386(clk,rst,matrix_A[386],matrix_B[186],mul_res1[386]);
multi_7x28 multi_7x28_mod_387(clk,rst,matrix_A[387],matrix_B[187],mul_res1[387]);
multi_7x28 multi_7x28_mod_388(clk,rst,matrix_A[388],matrix_B[188],mul_res1[388]);
multi_7x28 multi_7x28_mod_389(clk,rst,matrix_A[389],matrix_B[189],mul_res1[389]);
multi_7x28 multi_7x28_mod_390(clk,rst,matrix_A[390],matrix_B[190],mul_res1[390]);
multi_7x28 multi_7x28_mod_391(clk,rst,matrix_A[391],matrix_B[191],mul_res1[391]);
multi_7x28 multi_7x28_mod_392(clk,rst,matrix_A[392],matrix_B[192],mul_res1[392]);
multi_7x28 multi_7x28_mod_393(clk,rst,matrix_A[393],matrix_B[193],mul_res1[393]);
multi_7x28 multi_7x28_mod_394(clk,rst,matrix_A[394],matrix_B[194],mul_res1[394]);
multi_7x28 multi_7x28_mod_395(clk,rst,matrix_A[395],matrix_B[195],mul_res1[395]);
multi_7x28 multi_7x28_mod_396(clk,rst,matrix_A[396],matrix_B[196],mul_res1[396]);
multi_7x28 multi_7x28_mod_397(clk,rst,matrix_A[397],matrix_B[197],mul_res1[397]);
multi_7x28 multi_7x28_mod_398(clk,rst,matrix_A[398],matrix_B[198],mul_res1[398]);
multi_7x28 multi_7x28_mod_399(clk,rst,matrix_A[399],matrix_B[199],mul_res1[399]);
multi_7x28 multi_7x28_mod_400(clk,rst,matrix_A[400],matrix_B[0],mul_res1[400]);
multi_7x28 multi_7x28_mod_401(clk,rst,matrix_A[401],matrix_B[1],mul_res1[401]);
multi_7x28 multi_7x28_mod_402(clk,rst,matrix_A[402],matrix_B[2],mul_res1[402]);
multi_7x28 multi_7x28_mod_403(clk,rst,matrix_A[403],matrix_B[3],mul_res1[403]);
multi_7x28 multi_7x28_mod_404(clk,rst,matrix_A[404],matrix_B[4],mul_res1[404]);
multi_7x28 multi_7x28_mod_405(clk,rst,matrix_A[405],matrix_B[5],mul_res1[405]);
multi_7x28 multi_7x28_mod_406(clk,rst,matrix_A[406],matrix_B[6],mul_res1[406]);
multi_7x28 multi_7x28_mod_407(clk,rst,matrix_A[407],matrix_B[7],mul_res1[407]);
multi_7x28 multi_7x28_mod_408(clk,rst,matrix_A[408],matrix_B[8],mul_res1[408]);
multi_7x28 multi_7x28_mod_409(clk,rst,matrix_A[409],matrix_B[9],mul_res1[409]);
multi_7x28 multi_7x28_mod_410(clk,rst,matrix_A[410],matrix_B[10],mul_res1[410]);
multi_7x28 multi_7x28_mod_411(clk,rst,matrix_A[411],matrix_B[11],mul_res1[411]);
multi_7x28 multi_7x28_mod_412(clk,rst,matrix_A[412],matrix_B[12],mul_res1[412]);
multi_7x28 multi_7x28_mod_413(clk,rst,matrix_A[413],matrix_B[13],mul_res1[413]);
multi_7x28 multi_7x28_mod_414(clk,rst,matrix_A[414],matrix_B[14],mul_res1[414]);
multi_7x28 multi_7x28_mod_415(clk,rst,matrix_A[415],matrix_B[15],mul_res1[415]);
multi_7x28 multi_7x28_mod_416(clk,rst,matrix_A[416],matrix_B[16],mul_res1[416]);
multi_7x28 multi_7x28_mod_417(clk,rst,matrix_A[417],matrix_B[17],mul_res1[417]);
multi_7x28 multi_7x28_mod_418(clk,rst,matrix_A[418],matrix_B[18],mul_res1[418]);
multi_7x28 multi_7x28_mod_419(clk,rst,matrix_A[419],matrix_B[19],mul_res1[419]);
multi_7x28 multi_7x28_mod_420(clk,rst,matrix_A[420],matrix_B[20],mul_res1[420]);
multi_7x28 multi_7x28_mod_421(clk,rst,matrix_A[421],matrix_B[21],mul_res1[421]);
multi_7x28 multi_7x28_mod_422(clk,rst,matrix_A[422],matrix_B[22],mul_res1[422]);
multi_7x28 multi_7x28_mod_423(clk,rst,matrix_A[423],matrix_B[23],mul_res1[423]);
multi_7x28 multi_7x28_mod_424(clk,rst,matrix_A[424],matrix_B[24],mul_res1[424]);
multi_7x28 multi_7x28_mod_425(clk,rst,matrix_A[425],matrix_B[25],mul_res1[425]);
multi_7x28 multi_7x28_mod_426(clk,rst,matrix_A[426],matrix_B[26],mul_res1[426]);
multi_7x28 multi_7x28_mod_427(clk,rst,matrix_A[427],matrix_B[27],mul_res1[427]);
multi_7x28 multi_7x28_mod_428(clk,rst,matrix_A[428],matrix_B[28],mul_res1[428]);
multi_7x28 multi_7x28_mod_429(clk,rst,matrix_A[429],matrix_B[29],mul_res1[429]);
multi_7x28 multi_7x28_mod_430(clk,rst,matrix_A[430],matrix_B[30],mul_res1[430]);
multi_7x28 multi_7x28_mod_431(clk,rst,matrix_A[431],matrix_B[31],mul_res1[431]);
multi_7x28 multi_7x28_mod_432(clk,rst,matrix_A[432],matrix_B[32],mul_res1[432]);
multi_7x28 multi_7x28_mod_433(clk,rst,matrix_A[433],matrix_B[33],mul_res1[433]);
multi_7x28 multi_7x28_mod_434(clk,rst,matrix_A[434],matrix_B[34],mul_res1[434]);
multi_7x28 multi_7x28_mod_435(clk,rst,matrix_A[435],matrix_B[35],mul_res1[435]);
multi_7x28 multi_7x28_mod_436(clk,rst,matrix_A[436],matrix_B[36],mul_res1[436]);
multi_7x28 multi_7x28_mod_437(clk,rst,matrix_A[437],matrix_B[37],mul_res1[437]);
multi_7x28 multi_7x28_mod_438(clk,rst,matrix_A[438],matrix_B[38],mul_res1[438]);
multi_7x28 multi_7x28_mod_439(clk,rst,matrix_A[439],matrix_B[39],mul_res1[439]);
multi_7x28 multi_7x28_mod_440(clk,rst,matrix_A[440],matrix_B[40],mul_res1[440]);
multi_7x28 multi_7x28_mod_441(clk,rst,matrix_A[441],matrix_B[41],mul_res1[441]);
multi_7x28 multi_7x28_mod_442(clk,rst,matrix_A[442],matrix_B[42],mul_res1[442]);
multi_7x28 multi_7x28_mod_443(clk,rst,matrix_A[443],matrix_B[43],mul_res1[443]);
multi_7x28 multi_7x28_mod_444(clk,rst,matrix_A[444],matrix_B[44],mul_res1[444]);
multi_7x28 multi_7x28_mod_445(clk,rst,matrix_A[445],matrix_B[45],mul_res1[445]);
multi_7x28 multi_7x28_mod_446(clk,rst,matrix_A[446],matrix_B[46],mul_res1[446]);
multi_7x28 multi_7x28_mod_447(clk,rst,matrix_A[447],matrix_B[47],mul_res1[447]);
multi_7x28 multi_7x28_mod_448(clk,rst,matrix_A[448],matrix_B[48],mul_res1[448]);
multi_7x28 multi_7x28_mod_449(clk,rst,matrix_A[449],matrix_B[49],mul_res1[449]);
multi_7x28 multi_7x28_mod_450(clk,rst,matrix_A[450],matrix_B[50],mul_res1[450]);
multi_7x28 multi_7x28_mod_451(clk,rst,matrix_A[451],matrix_B[51],mul_res1[451]);
multi_7x28 multi_7x28_mod_452(clk,rst,matrix_A[452],matrix_B[52],mul_res1[452]);
multi_7x28 multi_7x28_mod_453(clk,rst,matrix_A[453],matrix_B[53],mul_res1[453]);
multi_7x28 multi_7x28_mod_454(clk,rst,matrix_A[454],matrix_B[54],mul_res1[454]);
multi_7x28 multi_7x28_mod_455(clk,rst,matrix_A[455],matrix_B[55],mul_res1[455]);
multi_7x28 multi_7x28_mod_456(clk,rst,matrix_A[456],matrix_B[56],mul_res1[456]);
multi_7x28 multi_7x28_mod_457(clk,rst,matrix_A[457],matrix_B[57],mul_res1[457]);
multi_7x28 multi_7x28_mod_458(clk,rst,matrix_A[458],matrix_B[58],mul_res1[458]);
multi_7x28 multi_7x28_mod_459(clk,rst,matrix_A[459],matrix_B[59],mul_res1[459]);
multi_7x28 multi_7x28_mod_460(clk,rst,matrix_A[460],matrix_B[60],mul_res1[460]);
multi_7x28 multi_7x28_mod_461(clk,rst,matrix_A[461],matrix_B[61],mul_res1[461]);
multi_7x28 multi_7x28_mod_462(clk,rst,matrix_A[462],matrix_B[62],mul_res1[462]);
multi_7x28 multi_7x28_mod_463(clk,rst,matrix_A[463],matrix_B[63],mul_res1[463]);
multi_7x28 multi_7x28_mod_464(clk,rst,matrix_A[464],matrix_B[64],mul_res1[464]);
multi_7x28 multi_7x28_mod_465(clk,rst,matrix_A[465],matrix_B[65],mul_res1[465]);
multi_7x28 multi_7x28_mod_466(clk,rst,matrix_A[466],matrix_B[66],mul_res1[466]);
multi_7x28 multi_7x28_mod_467(clk,rst,matrix_A[467],matrix_B[67],mul_res1[467]);
multi_7x28 multi_7x28_mod_468(clk,rst,matrix_A[468],matrix_B[68],mul_res1[468]);
multi_7x28 multi_7x28_mod_469(clk,rst,matrix_A[469],matrix_B[69],mul_res1[469]);
multi_7x28 multi_7x28_mod_470(clk,rst,matrix_A[470],matrix_B[70],mul_res1[470]);
multi_7x28 multi_7x28_mod_471(clk,rst,matrix_A[471],matrix_B[71],mul_res1[471]);
multi_7x28 multi_7x28_mod_472(clk,rst,matrix_A[472],matrix_B[72],mul_res1[472]);
multi_7x28 multi_7x28_mod_473(clk,rst,matrix_A[473],matrix_B[73],mul_res1[473]);
multi_7x28 multi_7x28_mod_474(clk,rst,matrix_A[474],matrix_B[74],mul_res1[474]);
multi_7x28 multi_7x28_mod_475(clk,rst,matrix_A[475],matrix_B[75],mul_res1[475]);
multi_7x28 multi_7x28_mod_476(clk,rst,matrix_A[476],matrix_B[76],mul_res1[476]);
multi_7x28 multi_7x28_mod_477(clk,rst,matrix_A[477],matrix_B[77],mul_res1[477]);
multi_7x28 multi_7x28_mod_478(clk,rst,matrix_A[478],matrix_B[78],mul_res1[478]);
multi_7x28 multi_7x28_mod_479(clk,rst,matrix_A[479],matrix_B[79],mul_res1[479]);
multi_7x28 multi_7x28_mod_480(clk,rst,matrix_A[480],matrix_B[80],mul_res1[480]);
multi_7x28 multi_7x28_mod_481(clk,rst,matrix_A[481],matrix_B[81],mul_res1[481]);
multi_7x28 multi_7x28_mod_482(clk,rst,matrix_A[482],matrix_B[82],mul_res1[482]);
multi_7x28 multi_7x28_mod_483(clk,rst,matrix_A[483],matrix_B[83],mul_res1[483]);
multi_7x28 multi_7x28_mod_484(clk,rst,matrix_A[484],matrix_B[84],mul_res1[484]);
multi_7x28 multi_7x28_mod_485(clk,rst,matrix_A[485],matrix_B[85],mul_res1[485]);
multi_7x28 multi_7x28_mod_486(clk,rst,matrix_A[486],matrix_B[86],mul_res1[486]);
multi_7x28 multi_7x28_mod_487(clk,rst,matrix_A[487],matrix_B[87],mul_res1[487]);
multi_7x28 multi_7x28_mod_488(clk,rst,matrix_A[488],matrix_B[88],mul_res1[488]);
multi_7x28 multi_7x28_mod_489(clk,rst,matrix_A[489],matrix_B[89],mul_res1[489]);
multi_7x28 multi_7x28_mod_490(clk,rst,matrix_A[490],matrix_B[90],mul_res1[490]);
multi_7x28 multi_7x28_mod_491(clk,rst,matrix_A[491],matrix_B[91],mul_res1[491]);
multi_7x28 multi_7x28_mod_492(clk,rst,matrix_A[492],matrix_B[92],mul_res1[492]);
multi_7x28 multi_7x28_mod_493(clk,rst,matrix_A[493],matrix_B[93],mul_res1[493]);
multi_7x28 multi_7x28_mod_494(clk,rst,matrix_A[494],matrix_B[94],mul_res1[494]);
multi_7x28 multi_7x28_mod_495(clk,rst,matrix_A[495],matrix_B[95],mul_res1[495]);
multi_7x28 multi_7x28_mod_496(clk,rst,matrix_A[496],matrix_B[96],mul_res1[496]);
multi_7x28 multi_7x28_mod_497(clk,rst,matrix_A[497],matrix_B[97],mul_res1[497]);
multi_7x28 multi_7x28_mod_498(clk,rst,matrix_A[498],matrix_B[98],mul_res1[498]);
multi_7x28 multi_7x28_mod_499(clk,rst,matrix_A[499],matrix_B[99],mul_res1[499]);
multi_7x28 multi_7x28_mod_500(clk,rst,matrix_A[500],matrix_B[100],mul_res1[500]);
multi_7x28 multi_7x28_mod_501(clk,rst,matrix_A[501],matrix_B[101],mul_res1[501]);
multi_7x28 multi_7x28_mod_502(clk,rst,matrix_A[502],matrix_B[102],mul_res1[502]);
multi_7x28 multi_7x28_mod_503(clk,rst,matrix_A[503],matrix_B[103],mul_res1[503]);
multi_7x28 multi_7x28_mod_504(clk,rst,matrix_A[504],matrix_B[104],mul_res1[504]);
multi_7x28 multi_7x28_mod_505(clk,rst,matrix_A[505],matrix_B[105],mul_res1[505]);
multi_7x28 multi_7x28_mod_506(clk,rst,matrix_A[506],matrix_B[106],mul_res1[506]);
multi_7x28 multi_7x28_mod_507(clk,rst,matrix_A[507],matrix_B[107],mul_res1[507]);
multi_7x28 multi_7x28_mod_508(clk,rst,matrix_A[508],matrix_B[108],mul_res1[508]);
multi_7x28 multi_7x28_mod_509(clk,rst,matrix_A[509],matrix_B[109],mul_res1[509]);
multi_7x28 multi_7x28_mod_510(clk,rst,matrix_A[510],matrix_B[110],mul_res1[510]);
multi_7x28 multi_7x28_mod_511(clk,rst,matrix_A[511],matrix_B[111],mul_res1[511]);
multi_7x28 multi_7x28_mod_512(clk,rst,matrix_A[512],matrix_B[112],mul_res1[512]);
multi_7x28 multi_7x28_mod_513(clk,rst,matrix_A[513],matrix_B[113],mul_res1[513]);
multi_7x28 multi_7x28_mod_514(clk,rst,matrix_A[514],matrix_B[114],mul_res1[514]);
multi_7x28 multi_7x28_mod_515(clk,rst,matrix_A[515],matrix_B[115],mul_res1[515]);
multi_7x28 multi_7x28_mod_516(clk,rst,matrix_A[516],matrix_B[116],mul_res1[516]);
multi_7x28 multi_7x28_mod_517(clk,rst,matrix_A[517],matrix_B[117],mul_res1[517]);
multi_7x28 multi_7x28_mod_518(clk,rst,matrix_A[518],matrix_B[118],mul_res1[518]);
multi_7x28 multi_7x28_mod_519(clk,rst,matrix_A[519],matrix_B[119],mul_res1[519]);
multi_7x28 multi_7x28_mod_520(clk,rst,matrix_A[520],matrix_B[120],mul_res1[520]);
multi_7x28 multi_7x28_mod_521(clk,rst,matrix_A[521],matrix_B[121],mul_res1[521]);
multi_7x28 multi_7x28_mod_522(clk,rst,matrix_A[522],matrix_B[122],mul_res1[522]);
multi_7x28 multi_7x28_mod_523(clk,rst,matrix_A[523],matrix_B[123],mul_res1[523]);
multi_7x28 multi_7x28_mod_524(clk,rst,matrix_A[524],matrix_B[124],mul_res1[524]);
multi_7x28 multi_7x28_mod_525(clk,rst,matrix_A[525],matrix_B[125],mul_res1[525]);
multi_7x28 multi_7x28_mod_526(clk,rst,matrix_A[526],matrix_B[126],mul_res1[526]);
multi_7x28 multi_7x28_mod_527(clk,rst,matrix_A[527],matrix_B[127],mul_res1[527]);
multi_7x28 multi_7x28_mod_528(clk,rst,matrix_A[528],matrix_B[128],mul_res1[528]);
multi_7x28 multi_7x28_mod_529(clk,rst,matrix_A[529],matrix_B[129],mul_res1[529]);
multi_7x28 multi_7x28_mod_530(clk,rst,matrix_A[530],matrix_B[130],mul_res1[530]);
multi_7x28 multi_7x28_mod_531(clk,rst,matrix_A[531],matrix_B[131],mul_res1[531]);
multi_7x28 multi_7x28_mod_532(clk,rst,matrix_A[532],matrix_B[132],mul_res1[532]);
multi_7x28 multi_7x28_mod_533(clk,rst,matrix_A[533],matrix_B[133],mul_res1[533]);
multi_7x28 multi_7x28_mod_534(clk,rst,matrix_A[534],matrix_B[134],mul_res1[534]);
multi_7x28 multi_7x28_mod_535(clk,rst,matrix_A[535],matrix_B[135],mul_res1[535]);
multi_7x28 multi_7x28_mod_536(clk,rst,matrix_A[536],matrix_B[136],mul_res1[536]);
multi_7x28 multi_7x28_mod_537(clk,rst,matrix_A[537],matrix_B[137],mul_res1[537]);
multi_7x28 multi_7x28_mod_538(clk,rst,matrix_A[538],matrix_B[138],mul_res1[538]);
multi_7x28 multi_7x28_mod_539(clk,rst,matrix_A[539],matrix_B[139],mul_res1[539]);
multi_7x28 multi_7x28_mod_540(clk,rst,matrix_A[540],matrix_B[140],mul_res1[540]);
multi_7x28 multi_7x28_mod_541(clk,rst,matrix_A[541],matrix_B[141],mul_res1[541]);
multi_7x28 multi_7x28_mod_542(clk,rst,matrix_A[542],matrix_B[142],mul_res1[542]);
multi_7x28 multi_7x28_mod_543(clk,rst,matrix_A[543],matrix_B[143],mul_res1[543]);
multi_7x28 multi_7x28_mod_544(clk,rst,matrix_A[544],matrix_B[144],mul_res1[544]);
multi_7x28 multi_7x28_mod_545(clk,rst,matrix_A[545],matrix_B[145],mul_res1[545]);
multi_7x28 multi_7x28_mod_546(clk,rst,matrix_A[546],matrix_B[146],mul_res1[546]);
multi_7x28 multi_7x28_mod_547(clk,rst,matrix_A[547],matrix_B[147],mul_res1[547]);
multi_7x28 multi_7x28_mod_548(clk,rst,matrix_A[548],matrix_B[148],mul_res1[548]);
multi_7x28 multi_7x28_mod_549(clk,rst,matrix_A[549],matrix_B[149],mul_res1[549]);
multi_7x28 multi_7x28_mod_550(clk,rst,matrix_A[550],matrix_B[150],mul_res1[550]);
multi_7x28 multi_7x28_mod_551(clk,rst,matrix_A[551],matrix_B[151],mul_res1[551]);
multi_7x28 multi_7x28_mod_552(clk,rst,matrix_A[552],matrix_B[152],mul_res1[552]);
multi_7x28 multi_7x28_mod_553(clk,rst,matrix_A[553],matrix_B[153],mul_res1[553]);
multi_7x28 multi_7x28_mod_554(clk,rst,matrix_A[554],matrix_B[154],mul_res1[554]);
multi_7x28 multi_7x28_mod_555(clk,rst,matrix_A[555],matrix_B[155],mul_res1[555]);
multi_7x28 multi_7x28_mod_556(clk,rst,matrix_A[556],matrix_B[156],mul_res1[556]);
multi_7x28 multi_7x28_mod_557(clk,rst,matrix_A[557],matrix_B[157],mul_res1[557]);
multi_7x28 multi_7x28_mod_558(clk,rst,matrix_A[558],matrix_B[158],mul_res1[558]);
multi_7x28 multi_7x28_mod_559(clk,rst,matrix_A[559],matrix_B[159],mul_res1[559]);
multi_7x28 multi_7x28_mod_560(clk,rst,matrix_A[560],matrix_B[160],mul_res1[560]);
multi_7x28 multi_7x28_mod_561(clk,rst,matrix_A[561],matrix_B[161],mul_res1[561]);
multi_7x28 multi_7x28_mod_562(clk,rst,matrix_A[562],matrix_B[162],mul_res1[562]);
multi_7x28 multi_7x28_mod_563(clk,rst,matrix_A[563],matrix_B[163],mul_res1[563]);
multi_7x28 multi_7x28_mod_564(clk,rst,matrix_A[564],matrix_B[164],mul_res1[564]);
multi_7x28 multi_7x28_mod_565(clk,rst,matrix_A[565],matrix_B[165],mul_res1[565]);
multi_7x28 multi_7x28_mod_566(clk,rst,matrix_A[566],matrix_B[166],mul_res1[566]);
multi_7x28 multi_7x28_mod_567(clk,rst,matrix_A[567],matrix_B[167],mul_res1[567]);
multi_7x28 multi_7x28_mod_568(clk,rst,matrix_A[568],matrix_B[168],mul_res1[568]);
multi_7x28 multi_7x28_mod_569(clk,rst,matrix_A[569],matrix_B[169],mul_res1[569]);
multi_7x28 multi_7x28_mod_570(clk,rst,matrix_A[570],matrix_B[170],mul_res1[570]);
multi_7x28 multi_7x28_mod_571(clk,rst,matrix_A[571],matrix_B[171],mul_res1[571]);
multi_7x28 multi_7x28_mod_572(clk,rst,matrix_A[572],matrix_B[172],mul_res1[572]);
multi_7x28 multi_7x28_mod_573(clk,rst,matrix_A[573],matrix_B[173],mul_res1[573]);
multi_7x28 multi_7x28_mod_574(clk,rst,matrix_A[574],matrix_B[174],mul_res1[574]);
multi_7x28 multi_7x28_mod_575(clk,rst,matrix_A[575],matrix_B[175],mul_res1[575]);
multi_7x28 multi_7x28_mod_576(clk,rst,matrix_A[576],matrix_B[176],mul_res1[576]);
multi_7x28 multi_7x28_mod_577(clk,rst,matrix_A[577],matrix_B[177],mul_res1[577]);
multi_7x28 multi_7x28_mod_578(clk,rst,matrix_A[578],matrix_B[178],mul_res1[578]);
multi_7x28 multi_7x28_mod_579(clk,rst,matrix_A[579],matrix_B[179],mul_res1[579]);
multi_7x28 multi_7x28_mod_580(clk,rst,matrix_A[580],matrix_B[180],mul_res1[580]);
multi_7x28 multi_7x28_mod_581(clk,rst,matrix_A[581],matrix_B[181],mul_res1[581]);
multi_7x28 multi_7x28_mod_582(clk,rst,matrix_A[582],matrix_B[182],mul_res1[582]);
multi_7x28 multi_7x28_mod_583(clk,rst,matrix_A[583],matrix_B[183],mul_res1[583]);
multi_7x28 multi_7x28_mod_584(clk,rst,matrix_A[584],matrix_B[184],mul_res1[584]);
multi_7x28 multi_7x28_mod_585(clk,rst,matrix_A[585],matrix_B[185],mul_res1[585]);
multi_7x28 multi_7x28_mod_586(clk,rst,matrix_A[586],matrix_B[186],mul_res1[586]);
multi_7x28 multi_7x28_mod_587(clk,rst,matrix_A[587],matrix_B[187],mul_res1[587]);
multi_7x28 multi_7x28_mod_588(clk,rst,matrix_A[588],matrix_B[188],mul_res1[588]);
multi_7x28 multi_7x28_mod_589(clk,rst,matrix_A[589],matrix_B[189],mul_res1[589]);
multi_7x28 multi_7x28_mod_590(clk,rst,matrix_A[590],matrix_B[190],mul_res1[590]);
multi_7x28 multi_7x28_mod_591(clk,rst,matrix_A[591],matrix_B[191],mul_res1[591]);
multi_7x28 multi_7x28_mod_592(clk,rst,matrix_A[592],matrix_B[192],mul_res1[592]);
multi_7x28 multi_7x28_mod_593(clk,rst,matrix_A[593],matrix_B[193],mul_res1[593]);
multi_7x28 multi_7x28_mod_594(clk,rst,matrix_A[594],matrix_B[194],mul_res1[594]);
multi_7x28 multi_7x28_mod_595(clk,rst,matrix_A[595],matrix_B[195],mul_res1[595]);
multi_7x28 multi_7x28_mod_596(clk,rst,matrix_A[596],matrix_B[196],mul_res1[596]);
multi_7x28 multi_7x28_mod_597(clk,rst,matrix_A[597],matrix_B[197],mul_res1[597]);
multi_7x28 multi_7x28_mod_598(clk,rst,matrix_A[598],matrix_B[198],mul_res1[598]);
multi_7x28 multi_7x28_mod_599(clk,rst,matrix_A[599],matrix_B[199],mul_res1[599]);
multi_7x28 multi_7x28_mod_600(clk,rst,matrix_A[600],matrix_B[0],mul_res1[600]);
multi_7x28 multi_7x28_mod_601(clk,rst,matrix_A[601],matrix_B[1],mul_res1[601]);
multi_7x28 multi_7x28_mod_602(clk,rst,matrix_A[602],matrix_B[2],mul_res1[602]);
multi_7x28 multi_7x28_mod_603(clk,rst,matrix_A[603],matrix_B[3],mul_res1[603]);
multi_7x28 multi_7x28_mod_604(clk,rst,matrix_A[604],matrix_B[4],mul_res1[604]);
multi_7x28 multi_7x28_mod_605(clk,rst,matrix_A[605],matrix_B[5],mul_res1[605]);
multi_7x28 multi_7x28_mod_606(clk,rst,matrix_A[606],matrix_B[6],mul_res1[606]);
multi_7x28 multi_7x28_mod_607(clk,rst,matrix_A[607],matrix_B[7],mul_res1[607]);
multi_7x28 multi_7x28_mod_608(clk,rst,matrix_A[608],matrix_B[8],mul_res1[608]);
multi_7x28 multi_7x28_mod_609(clk,rst,matrix_A[609],matrix_B[9],mul_res1[609]);
multi_7x28 multi_7x28_mod_610(clk,rst,matrix_A[610],matrix_B[10],mul_res1[610]);
multi_7x28 multi_7x28_mod_611(clk,rst,matrix_A[611],matrix_B[11],mul_res1[611]);
multi_7x28 multi_7x28_mod_612(clk,rst,matrix_A[612],matrix_B[12],mul_res1[612]);
multi_7x28 multi_7x28_mod_613(clk,rst,matrix_A[613],matrix_B[13],mul_res1[613]);
multi_7x28 multi_7x28_mod_614(clk,rst,matrix_A[614],matrix_B[14],mul_res1[614]);
multi_7x28 multi_7x28_mod_615(clk,rst,matrix_A[615],matrix_B[15],mul_res1[615]);
multi_7x28 multi_7x28_mod_616(clk,rst,matrix_A[616],matrix_B[16],mul_res1[616]);
multi_7x28 multi_7x28_mod_617(clk,rst,matrix_A[617],matrix_B[17],mul_res1[617]);
multi_7x28 multi_7x28_mod_618(clk,rst,matrix_A[618],matrix_B[18],mul_res1[618]);
multi_7x28 multi_7x28_mod_619(clk,rst,matrix_A[619],matrix_B[19],mul_res1[619]);
multi_7x28 multi_7x28_mod_620(clk,rst,matrix_A[620],matrix_B[20],mul_res1[620]);
multi_7x28 multi_7x28_mod_621(clk,rst,matrix_A[621],matrix_B[21],mul_res1[621]);
multi_7x28 multi_7x28_mod_622(clk,rst,matrix_A[622],matrix_B[22],mul_res1[622]);
multi_7x28 multi_7x28_mod_623(clk,rst,matrix_A[623],matrix_B[23],mul_res1[623]);
multi_7x28 multi_7x28_mod_624(clk,rst,matrix_A[624],matrix_B[24],mul_res1[624]);
multi_7x28 multi_7x28_mod_625(clk,rst,matrix_A[625],matrix_B[25],mul_res1[625]);
multi_7x28 multi_7x28_mod_626(clk,rst,matrix_A[626],matrix_B[26],mul_res1[626]);
multi_7x28 multi_7x28_mod_627(clk,rst,matrix_A[627],matrix_B[27],mul_res1[627]);
multi_7x28 multi_7x28_mod_628(clk,rst,matrix_A[628],matrix_B[28],mul_res1[628]);
multi_7x28 multi_7x28_mod_629(clk,rst,matrix_A[629],matrix_B[29],mul_res1[629]);
multi_7x28 multi_7x28_mod_630(clk,rst,matrix_A[630],matrix_B[30],mul_res1[630]);
multi_7x28 multi_7x28_mod_631(clk,rst,matrix_A[631],matrix_B[31],mul_res1[631]);
multi_7x28 multi_7x28_mod_632(clk,rst,matrix_A[632],matrix_B[32],mul_res1[632]);
multi_7x28 multi_7x28_mod_633(clk,rst,matrix_A[633],matrix_B[33],mul_res1[633]);
multi_7x28 multi_7x28_mod_634(clk,rst,matrix_A[634],matrix_B[34],mul_res1[634]);
multi_7x28 multi_7x28_mod_635(clk,rst,matrix_A[635],matrix_B[35],mul_res1[635]);
multi_7x28 multi_7x28_mod_636(clk,rst,matrix_A[636],matrix_B[36],mul_res1[636]);
multi_7x28 multi_7x28_mod_637(clk,rst,matrix_A[637],matrix_B[37],mul_res1[637]);
multi_7x28 multi_7x28_mod_638(clk,rst,matrix_A[638],matrix_B[38],mul_res1[638]);
multi_7x28 multi_7x28_mod_639(clk,rst,matrix_A[639],matrix_B[39],mul_res1[639]);
multi_7x28 multi_7x28_mod_640(clk,rst,matrix_A[640],matrix_B[40],mul_res1[640]);
multi_7x28 multi_7x28_mod_641(clk,rst,matrix_A[641],matrix_B[41],mul_res1[641]);
multi_7x28 multi_7x28_mod_642(clk,rst,matrix_A[642],matrix_B[42],mul_res1[642]);
multi_7x28 multi_7x28_mod_643(clk,rst,matrix_A[643],matrix_B[43],mul_res1[643]);
multi_7x28 multi_7x28_mod_644(clk,rst,matrix_A[644],matrix_B[44],mul_res1[644]);
multi_7x28 multi_7x28_mod_645(clk,rst,matrix_A[645],matrix_B[45],mul_res1[645]);
multi_7x28 multi_7x28_mod_646(clk,rst,matrix_A[646],matrix_B[46],mul_res1[646]);
multi_7x28 multi_7x28_mod_647(clk,rst,matrix_A[647],matrix_B[47],mul_res1[647]);
multi_7x28 multi_7x28_mod_648(clk,rst,matrix_A[648],matrix_B[48],mul_res1[648]);
multi_7x28 multi_7x28_mod_649(clk,rst,matrix_A[649],matrix_B[49],mul_res1[649]);
multi_7x28 multi_7x28_mod_650(clk,rst,matrix_A[650],matrix_B[50],mul_res1[650]);
multi_7x28 multi_7x28_mod_651(clk,rst,matrix_A[651],matrix_B[51],mul_res1[651]);
multi_7x28 multi_7x28_mod_652(clk,rst,matrix_A[652],matrix_B[52],mul_res1[652]);
multi_7x28 multi_7x28_mod_653(clk,rst,matrix_A[653],matrix_B[53],mul_res1[653]);
multi_7x28 multi_7x28_mod_654(clk,rst,matrix_A[654],matrix_B[54],mul_res1[654]);
multi_7x28 multi_7x28_mod_655(clk,rst,matrix_A[655],matrix_B[55],mul_res1[655]);
multi_7x28 multi_7x28_mod_656(clk,rst,matrix_A[656],matrix_B[56],mul_res1[656]);
multi_7x28 multi_7x28_mod_657(clk,rst,matrix_A[657],matrix_B[57],mul_res1[657]);
multi_7x28 multi_7x28_mod_658(clk,rst,matrix_A[658],matrix_B[58],mul_res1[658]);
multi_7x28 multi_7x28_mod_659(clk,rst,matrix_A[659],matrix_B[59],mul_res1[659]);
multi_7x28 multi_7x28_mod_660(clk,rst,matrix_A[660],matrix_B[60],mul_res1[660]);
multi_7x28 multi_7x28_mod_661(clk,rst,matrix_A[661],matrix_B[61],mul_res1[661]);
multi_7x28 multi_7x28_mod_662(clk,rst,matrix_A[662],matrix_B[62],mul_res1[662]);
multi_7x28 multi_7x28_mod_663(clk,rst,matrix_A[663],matrix_B[63],mul_res1[663]);
multi_7x28 multi_7x28_mod_664(clk,rst,matrix_A[664],matrix_B[64],mul_res1[664]);
multi_7x28 multi_7x28_mod_665(clk,rst,matrix_A[665],matrix_B[65],mul_res1[665]);
multi_7x28 multi_7x28_mod_666(clk,rst,matrix_A[666],matrix_B[66],mul_res1[666]);
multi_7x28 multi_7x28_mod_667(clk,rst,matrix_A[667],matrix_B[67],mul_res1[667]);
multi_7x28 multi_7x28_mod_668(clk,rst,matrix_A[668],matrix_B[68],mul_res1[668]);
multi_7x28 multi_7x28_mod_669(clk,rst,matrix_A[669],matrix_B[69],mul_res1[669]);
multi_7x28 multi_7x28_mod_670(clk,rst,matrix_A[670],matrix_B[70],mul_res1[670]);
multi_7x28 multi_7x28_mod_671(clk,rst,matrix_A[671],matrix_B[71],mul_res1[671]);
multi_7x28 multi_7x28_mod_672(clk,rst,matrix_A[672],matrix_B[72],mul_res1[672]);
multi_7x28 multi_7x28_mod_673(clk,rst,matrix_A[673],matrix_B[73],mul_res1[673]);
multi_7x28 multi_7x28_mod_674(clk,rst,matrix_A[674],matrix_B[74],mul_res1[674]);
multi_7x28 multi_7x28_mod_675(clk,rst,matrix_A[675],matrix_B[75],mul_res1[675]);
multi_7x28 multi_7x28_mod_676(clk,rst,matrix_A[676],matrix_B[76],mul_res1[676]);
multi_7x28 multi_7x28_mod_677(clk,rst,matrix_A[677],matrix_B[77],mul_res1[677]);
multi_7x28 multi_7x28_mod_678(clk,rst,matrix_A[678],matrix_B[78],mul_res1[678]);
multi_7x28 multi_7x28_mod_679(clk,rst,matrix_A[679],matrix_B[79],mul_res1[679]);
multi_7x28 multi_7x28_mod_680(clk,rst,matrix_A[680],matrix_B[80],mul_res1[680]);
multi_7x28 multi_7x28_mod_681(clk,rst,matrix_A[681],matrix_B[81],mul_res1[681]);
multi_7x28 multi_7x28_mod_682(clk,rst,matrix_A[682],matrix_B[82],mul_res1[682]);
multi_7x28 multi_7x28_mod_683(clk,rst,matrix_A[683],matrix_B[83],mul_res1[683]);
multi_7x28 multi_7x28_mod_684(clk,rst,matrix_A[684],matrix_B[84],mul_res1[684]);
multi_7x28 multi_7x28_mod_685(clk,rst,matrix_A[685],matrix_B[85],mul_res1[685]);
multi_7x28 multi_7x28_mod_686(clk,rst,matrix_A[686],matrix_B[86],mul_res1[686]);
multi_7x28 multi_7x28_mod_687(clk,rst,matrix_A[687],matrix_B[87],mul_res1[687]);
multi_7x28 multi_7x28_mod_688(clk,rst,matrix_A[688],matrix_B[88],mul_res1[688]);
multi_7x28 multi_7x28_mod_689(clk,rst,matrix_A[689],matrix_B[89],mul_res1[689]);
multi_7x28 multi_7x28_mod_690(clk,rst,matrix_A[690],matrix_B[90],mul_res1[690]);
multi_7x28 multi_7x28_mod_691(clk,rst,matrix_A[691],matrix_B[91],mul_res1[691]);
multi_7x28 multi_7x28_mod_692(clk,rst,matrix_A[692],matrix_B[92],mul_res1[692]);
multi_7x28 multi_7x28_mod_693(clk,rst,matrix_A[693],matrix_B[93],mul_res1[693]);
multi_7x28 multi_7x28_mod_694(clk,rst,matrix_A[694],matrix_B[94],mul_res1[694]);
multi_7x28 multi_7x28_mod_695(clk,rst,matrix_A[695],matrix_B[95],mul_res1[695]);
multi_7x28 multi_7x28_mod_696(clk,rst,matrix_A[696],matrix_B[96],mul_res1[696]);
multi_7x28 multi_7x28_mod_697(clk,rst,matrix_A[697],matrix_B[97],mul_res1[697]);
multi_7x28 multi_7x28_mod_698(clk,rst,matrix_A[698],matrix_B[98],mul_res1[698]);
multi_7x28 multi_7x28_mod_699(clk,rst,matrix_A[699],matrix_B[99],mul_res1[699]);
multi_7x28 multi_7x28_mod_700(clk,rst,matrix_A[700],matrix_B[100],mul_res1[700]);
multi_7x28 multi_7x28_mod_701(clk,rst,matrix_A[701],matrix_B[101],mul_res1[701]);
multi_7x28 multi_7x28_mod_702(clk,rst,matrix_A[702],matrix_B[102],mul_res1[702]);
multi_7x28 multi_7x28_mod_703(clk,rst,matrix_A[703],matrix_B[103],mul_res1[703]);
multi_7x28 multi_7x28_mod_704(clk,rst,matrix_A[704],matrix_B[104],mul_res1[704]);
multi_7x28 multi_7x28_mod_705(clk,rst,matrix_A[705],matrix_B[105],mul_res1[705]);
multi_7x28 multi_7x28_mod_706(clk,rst,matrix_A[706],matrix_B[106],mul_res1[706]);
multi_7x28 multi_7x28_mod_707(clk,rst,matrix_A[707],matrix_B[107],mul_res1[707]);
multi_7x28 multi_7x28_mod_708(clk,rst,matrix_A[708],matrix_B[108],mul_res1[708]);
multi_7x28 multi_7x28_mod_709(clk,rst,matrix_A[709],matrix_B[109],mul_res1[709]);
multi_7x28 multi_7x28_mod_710(clk,rst,matrix_A[710],matrix_B[110],mul_res1[710]);
multi_7x28 multi_7x28_mod_711(clk,rst,matrix_A[711],matrix_B[111],mul_res1[711]);
multi_7x28 multi_7x28_mod_712(clk,rst,matrix_A[712],matrix_B[112],mul_res1[712]);
multi_7x28 multi_7x28_mod_713(clk,rst,matrix_A[713],matrix_B[113],mul_res1[713]);
multi_7x28 multi_7x28_mod_714(clk,rst,matrix_A[714],matrix_B[114],mul_res1[714]);
multi_7x28 multi_7x28_mod_715(clk,rst,matrix_A[715],matrix_B[115],mul_res1[715]);
multi_7x28 multi_7x28_mod_716(clk,rst,matrix_A[716],matrix_B[116],mul_res1[716]);
multi_7x28 multi_7x28_mod_717(clk,rst,matrix_A[717],matrix_B[117],mul_res1[717]);
multi_7x28 multi_7x28_mod_718(clk,rst,matrix_A[718],matrix_B[118],mul_res1[718]);
multi_7x28 multi_7x28_mod_719(clk,rst,matrix_A[719],matrix_B[119],mul_res1[719]);
multi_7x28 multi_7x28_mod_720(clk,rst,matrix_A[720],matrix_B[120],mul_res1[720]);
multi_7x28 multi_7x28_mod_721(clk,rst,matrix_A[721],matrix_B[121],mul_res1[721]);
multi_7x28 multi_7x28_mod_722(clk,rst,matrix_A[722],matrix_B[122],mul_res1[722]);
multi_7x28 multi_7x28_mod_723(clk,rst,matrix_A[723],matrix_B[123],mul_res1[723]);
multi_7x28 multi_7x28_mod_724(clk,rst,matrix_A[724],matrix_B[124],mul_res1[724]);
multi_7x28 multi_7x28_mod_725(clk,rst,matrix_A[725],matrix_B[125],mul_res1[725]);
multi_7x28 multi_7x28_mod_726(clk,rst,matrix_A[726],matrix_B[126],mul_res1[726]);
multi_7x28 multi_7x28_mod_727(clk,rst,matrix_A[727],matrix_B[127],mul_res1[727]);
multi_7x28 multi_7x28_mod_728(clk,rst,matrix_A[728],matrix_B[128],mul_res1[728]);
multi_7x28 multi_7x28_mod_729(clk,rst,matrix_A[729],matrix_B[129],mul_res1[729]);
multi_7x28 multi_7x28_mod_730(clk,rst,matrix_A[730],matrix_B[130],mul_res1[730]);
multi_7x28 multi_7x28_mod_731(clk,rst,matrix_A[731],matrix_B[131],mul_res1[731]);
multi_7x28 multi_7x28_mod_732(clk,rst,matrix_A[732],matrix_B[132],mul_res1[732]);
multi_7x28 multi_7x28_mod_733(clk,rst,matrix_A[733],matrix_B[133],mul_res1[733]);
multi_7x28 multi_7x28_mod_734(clk,rst,matrix_A[734],matrix_B[134],mul_res1[734]);
multi_7x28 multi_7x28_mod_735(clk,rst,matrix_A[735],matrix_B[135],mul_res1[735]);
multi_7x28 multi_7x28_mod_736(clk,rst,matrix_A[736],matrix_B[136],mul_res1[736]);
multi_7x28 multi_7x28_mod_737(clk,rst,matrix_A[737],matrix_B[137],mul_res1[737]);
multi_7x28 multi_7x28_mod_738(clk,rst,matrix_A[738],matrix_B[138],mul_res1[738]);
multi_7x28 multi_7x28_mod_739(clk,rst,matrix_A[739],matrix_B[139],mul_res1[739]);
multi_7x28 multi_7x28_mod_740(clk,rst,matrix_A[740],matrix_B[140],mul_res1[740]);
multi_7x28 multi_7x28_mod_741(clk,rst,matrix_A[741],matrix_B[141],mul_res1[741]);
multi_7x28 multi_7x28_mod_742(clk,rst,matrix_A[742],matrix_B[142],mul_res1[742]);
multi_7x28 multi_7x28_mod_743(clk,rst,matrix_A[743],matrix_B[143],mul_res1[743]);
multi_7x28 multi_7x28_mod_744(clk,rst,matrix_A[744],matrix_B[144],mul_res1[744]);
multi_7x28 multi_7x28_mod_745(clk,rst,matrix_A[745],matrix_B[145],mul_res1[745]);
multi_7x28 multi_7x28_mod_746(clk,rst,matrix_A[746],matrix_B[146],mul_res1[746]);
multi_7x28 multi_7x28_mod_747(clk,rst,matrix_A[747],matrix_B[147],mul_res1[747]);
multi_7x28 multi_7x28_mod_748(clk,rst,matrix_A[748],matrix_B[148],mul_res1[748]);
multi_7x28 multi_7x28_mod_749(clk,rst,matrix_A[749],matrix_B[149],mul_res1[749]);
multi_7x28 multi_7x28_mod_750(clk,rst,matrix_A[750],matrix_B[150],mul_res1[750]);
multi_7x28 multi_7x28_mod_751(clk,rst,matrix_A[751],matrix_B[151],mul_res1[751]);
multi_7x28 multi_7x28_mod_752(clk,rst,matrix_A[752],matrix_B[152],mul_res1[752]);
multi_7x28 multi_7x28_mod_753(clk,rst,matrix_A[753],matrix_B[153],mul_res1[753]);
multi_7x28 multi_7x28_mod_754(clk,rst,matrix_A[754],matrix_B[154],mul_res1[754]);
multi_7x28 multi_7x28_mod_755(clk,rst,matrix_A[755],matrix_B[155],mul_res1[755]);
multi_7x28 multi_7x28_mod_756(clk,rst,matrix_A[756],matrix_B[156],mul_res1[756]);
multi_7x28 multi_7x28_mod_757(clk,rst,matrix_A[757],matrix_B[157],mul_res1[757]);
multi_7x28 multi_7x28_mod_758(clk,rst,matrix_A[758],matrix_B[158],mul_res1[758]);
multi_7x28 multi_7x28_mod_759(clk,rst,matrix_A[759],matrix_B[159],mul_res1[759]);
multi_7x28 multi_7x28_mod_760(clk,rst,matrix_A[760],matrix_B[160],mul_res1[760]);
multi_7x28 multi_7x28_mod_761(clk,rst,matrix_A[761],matrix_B[161],mul_res1[761]);
multi_7x28 multi_7x28_mod_762(clk,rst,matrix_A[762],matrix_B[162],mul_res1[762]);
multi_7x28 multi_7x28_mod_763(clk,rst,matrix_A[763],matrix_B[163],mul_res1[763]);
multi_7x28 multi_7x28_mod_764(clk,rst,matrix_A[764],matrix_B[164],mul_res1[764]);
multi_7x28 multi_7x28_mod_765(clk,rst,matrix_A[765],matrix_B[165],mul_res1[765]);
multi_7x28 multi_7x28_mod_766(clk,rst,matrix_A[766],matrix_B[166],mul_res1[766]);
multi_7x28 multi_7x28_mod_767(clk,rst,matrix_A[767],matrix_B[167],mul_res1[767]);
multi_7x28 multi_7x28_mod_768(clk,rst,matrix_A[768],matrix_B[168],mul_res1[768]);
multi_7x28 multi_7x28_mod_769(clk,rst,matrix_A[769],matrix_B[169],mul_res1[769]);
multi_7x28 multi_7x28_mod_770(clk,rst,matrix_A[770],matrix_B[170],mul_res1[770]);
multi_7x28 multi_7x28_mod_771(clk,rst,matrix_A[771],matrix_B[171],mul_res1[771]);
multi_7x28 multi_7x28_mod_772(clk,rst,matrix_A[772],matrix_B[172],mul_res1[772]);
multi_7x28 multi_7x28_mod_773(clk,rst,matrix_A[773],matrix_B[173],mul_res1[773]);
multi_7x28 multi_7x28_mod_774(clk,rst,matrix_A[774],matrix_B[174],mul_res1[774]);
multi_7x28 multi_7x28_mod_775(clk,rst,matrix_A[775],matrix_B[175],mul_res1[775]);
multi_7x28 multi_7x28_mod_776(clk,rst,matrix_A[776],matrix_B[176],mul_res1[776]);
multi_7x28 multi_7x28_mod_777(clk,rst,matrix_A[777],matrix_B[177],mul_res1[777]);
multi_7x28 multi_7x28_mod_778(clk,rst,matrix_A[778],matrix_B[178],mul_res1[778]);
multi_7x28 multi_7x28_mod_779(clk,rst,matrix_A[779],matrix_B[179],mul_res1[779]);
multi_7x28 multi_7x28_mod_780(clk,rst,matrix_A[780],matrix_B[180],mul_res1[780]);
multi_7x28 multi_7x28_mod_781(clk,rst,matrix_A[781],matrix_B[181],mul_res1[781]);
multi_7x28 multi_7x28_mod_782(clk,rst,matrix_A[782],matrix_B[182],mul_res1[782]);
multi_7x28 multi_7x28_mod_783(clk,rst,matrix_A[783],matrix_B[183],mul_res1[783]);
multi_7x28 multi_7x28_mod_784(clk,rst,matrix_A[784],matrix_B[184],mul_res1[784]);
multi_7x28 multi_7x28_mod_785(clk,rst,matrix_A[785],matrix_B[185],mul_res1[785]);
multi_7x28 multi_7x28_mod_786(clk,rst,matrix_A[786],matrix_B[186],mul_res1[786]);
multi_7x28 multi_7x28_mod_787(clk,rst,matrix_A[787],matrix_B[187],mul_res1[787]);
multi_7x28 multi_7x28_mod_788(clk,rst,matrix_A[788],matrix_B[188],mul_res1[788]);
multi_7x28 multi_7x28_mod_789(clk,rst,matrix_A[789],matrix_B[189],mul_res1[789]);
multi_7x28 multi_7x28_mod_790(clk,rst,matrix_A[790],matrix_B[190],mul_res1[790]);
multi_7x28 multi_7x28_mod_791(clk,rst,matrix_A[791],matrix_B[191],mul_res1[791]);
multi_7x28 multi_7x28_mod_792(clk,rst,matrix_A[792],matrix_B[192],mul_res1[792]);
multi_7x28 multi_7x28_mod_793(clk,rst,matrix_A[793],matrix_B[193],mul_res1[793]);
multi_7x28 multi_7x28_mod_794(clk,rst,matrix_A[794],matrix_B[194],mul_res1[794]);
multi_7x28 multi_7x28_mod_795(clk,rst,matrix_A[795],matrix_B[195],mul_res1[795]);
multi_7x28 multi_7x28_mod_796(clk,rst,matrix_A[796],matrix_B[196],mul_res1[796]);
multi_7x28 multi_7x28_mod_797(clk,rst,matrix_A[797],matrix_B[197],mul_res1[797]);
multi_7x28 multi_7x28_mod_798(clk,rst,matrix_A[798],matrix_B[198],mul_res1[798]);
multi_7x28 multi_7x28_mod_799(clk,rst,matrix_A[799],matrix_B[199],mul_res1[799]);
multi_7x28 multi_7x28_mod_800(clk,rst,matrix_A[800],matrix_B[0],mul_res1[800]);
multi_7x28 multi_7x28_mod_801(clk,rst,matrix_A[801],matrix_B[1],mul_res1[801]);
multi_7x28 multi_7x28_mod_802(clk,rst,matrix_A[802],matrix_B[2],mul_res1[802]);
multi_7x28 multi_7x28_mod_803(clk,rst,matrix_A[803],matrix_B[3],mul_res1[803]);
multi_7x28 multi_7x28_mod_804(clk,rst,matrix_A[804],matrix_B[4],mul_res1[804]);
multi_7x28 multi_7x28_mod_805(clk,rst,matrix_A[805],matrix_B[5],mul_res1[805]);
multi_7x28 multi_7x28_mod_806(clk,rst,matrix_A[806],matrix_B[6],mul_res1[806]);
multi_7x28 multi_7x28_mod_807(clk,rst,matrix_A[807],matrix_B[7],mul_res1[807]);
multi_7x28 multi_7x28_mod_808(clk,rst,matrix_A[808],matrix_B[8],mul_res1[808]);
multi_7x28 multi_7x28_mod_809(clk,rst,matrix_A[809],matrix_B[9],mul_res1[809]);
multi_7x28 multi_7x28_mod_810(clk,rst,matrix_A[810],matrix_B[10],mul_res1[810]);
multi_7x28 multi_7x28_mod_811(clk,rst,matrix_A[811],matrix_B[11],mul_res1[811]);
multi_7x28 multi_7x28_mod_812(clk,rst,matrix_A[812],matrix_B[12],mul_res1[812]);
multi_7x28 multi_7x28_mod_813(clk,rst,matrix_A[813],matrix_B[13],mul_res1[813]);
multi_7x28 multi_7x28_mod_814(clk,rst,matrix_A[814],matrix_B[14],mul_res1[814]);
multi_7x28 multi_7x28_mod_815(clk,rst,matrix_A[815],matrix_B[15],mul_res1[815]);
multi_7x28 multi_7x28_mod_816(clk,rst,matrix_A[816],matrix_B[16],mul_res1[816]);
multi_7x28 multi_7x28_mod_817(clk,rst,matrix_A[817],matrix_B[17],mul_res1[817]);
multi_7x28 multi_7x28_mod_818(clk,rst,matrix_A[818],matrix_B[18],mul_res1[818]);
multi_7x28 multi_7x28_mod_819(clk,rst,matrix_A[819],matrix_B[19],mul_res1[819]);
multi_7x28 multi_7x28_mod_820(clk,rst,matrix_A[820],matrix_B[20],mul_res1[820]);
multi_7x28 multi_7x28_mod_821(clk,rst,matrix_A[821],matrix_B[21],mul_res1[821]);
multi_7x28 multi_7x28_mod_822(clk,rst,matrix_A[822],matrix_B[22],mul_res1[822]);
multi_7x28 multi_7x28_mod_823(clk,rst,matrix_A[823],matrix_B[23],mul_res1[823]);
multi_7x28 multi_7x28_mod_824(clk,rst,matrix_A[824],matrix_B[24],mul_res1[824]);
multi_7x28 multi_7x28_mod_825(clk,rst,matrix_A[825],matrix_B[25],mul_res1[825]);
multi_7x28 multi_7x28_mod_826(clk,rst,matrix_A[826],matrix_B[26],mul_res1[826]);
multi_7x28 multi_7x28_mod_827(clk,rst,matrix_A[827],matrix_B[27],mul_res1[827]);
multi_7x28 multi_7x28_mod_828(clk,rst,matrix_A[828],matrix_B[28],mul_res1[828]);
multi_7x28 multi_7x28_mod_829(clk,rst,matrix_A[829],matrix_B[29],mul_res1[829]);
multi_7x28 multi_7x28_mod_830(clk,rst,matrix_A[830],matrix_B[30],mul_res1[830]);
multi_7x28 multi_7x28_mod_831(clk,rst,matrix_A[831],matrix_B[31],mul_res1[831]);
multi_7x28 multi_7x28_mod_832(clk,rst,matrix_A[832],matrix_B[32],mul_res1[832]);
multi_7x28 multi_7x28_mod_833(clk,rst,matrix_A[833],matrix_B[33],mul_res1[833]);
multi_7x28 multi_7x28_mod_834(clk,rst,matrix_A[834],matrix_B[34],mul_res1[834]);
multi_7x28 multi_7x28_mod_835(clk,rst,matrix_A[835],matrix_B[35],mul_res1[835]);
multi_7x28 multi_7x28_mod_836(clk,rst,matrix_A[836],matrix_B[36],mul_res1[836]);
multi_7x28 multi_7x28_mod_837(clk,rst,matrix_A[837],matrix_B[37],mul_res1[837]);
multi_7x28 multi_7x28_mod_838(clk,rst,matrix_A[838],matrix_B[38],mul_res1[838]);
multi_7x28 multi_7x28_mod_839(clk,rst,matrix_A[839],matrix_B[39],mul_res1[839]);
multi_7x28 multi_7x28_mod_840(clk,rst,matrix_A[840],matrix_B[40],mul_res1[840]);
multi_7x28 multi_7x28_mod_841(clk,rst,matrix_A[841],matrix_B[41],mul_res1[841]);
multi_7x28 multi_7x28_mod_842(clk,rst,matrix_A[842],matrix_B[42],mul_res1[842]);
multi_7x28 multi_7x28_mod_843(clk,rst,matrix_A[843],matrix_B[43],mul_res1[843]);
multi_7x28 multi_7x28_mod_844(clk,rst,matrix_A[844],matrix_B[44],mul_res1[844]);
multi_7x28 multi_7x28_mod_845(clk,rst,matrix_A[845],matrix_B[45],mul_res1[845]);
multi_7x28 multi_7x28_mod_846(clk,rst,matrix_A[846],matrix_B[46],mul_res1[846]);
multi_7x28 multi_7x28_mod_847(clk,rst,matrix_A[847],matrix_B[47],mul_res1[847]);
multi_7x28 multi_7x28_mod_848(clk,rst,matrix_A[848],matrix_B[48],mul_res1[848]);
multi_7x28 multi_7x28_mod_849(clk,rst,matrix_A[849],matrix_B[49],mul_res1[849]);
multi_7x28 multi_7x28_mod_850(clk,rst,matrix_A[850],matrix_B[50],mul_res1[850]);
multi_7x28 multi_7x28_mod_851(clk,rst,matrix_A[851],matrix_B[51],mul_res1[851]);
multi_7x28 multi_7x28_mod_852(clk,rst,matrix_A[852],matrix_B[52],mul_res1[852]);
multi_7x28 multi_7x28_mod_853(clk,rst,matrix_A[853],matrix_B[53],mul_res1[853]);
multi_7x28 multi_7x28_mod_854(clk,rst,matrix_A[854],matrix_B[54],mul_res1[854]);
multi_7x28 multi_7x28_mod_855(clk,rst,matrix_A[855],matrix_B[55],mul_res1[855]);
multi_7x28 multi_7x28_mod_856(clk,rst,matrix_A[856],matrix_B[56],mul_res1[856]);
multi_7x28 multi_7x28_mod_857(clk,rst,matrix_A[857],matrix_B[57],mul_res1[857]);
multi_7x28 multi_7x28_mod_858(clk,rst,matrix_A[858],matrix_B[58],mul_res1[858]);
multi_7x28 multi_7x28_mod_859(clk,rst,matrix_A[859],matrix_B[59],mul_res1[859]);
multi_7x28 multi_7x28_mod_860(clk,rst,matrix_A[860],matrix_B[60],mul_res1[860]);
multi_7x28 multi_7x28_mod_861(clk,rst,matrix_A[861],matrix_B[61],mul_res1[861]);
multi_7x28 multi_7x28_mod_862(clk,rst,matrix_A[862],matrix_B[62],mul_res1[862]);
multi_7x28 multi_7x28_mod_863(clk,rst,matrix_A[863],matrix_B[63],mul_res1[863]);
multi_7x28 multi_7x28_mod_864(clk,rst,matrix_A[864],matrix_B[64],mul_res1[864]);
multi_7x28 multi_7x28_mod_865(clk,rst,matrix_A[865],matrix_B[65],mul_res1[865]);
multi_7x28 multi_7x28_mod_866(clk,rst,matrix_A[866],matrix_B[66],mul_res1[866]);
multi_7x28 multi_7x28_mod_867(clk,rst,matrix_A[867],matrix_B[67],mul_res1[867]);
multi_7x28 multi_7x28_mod_868(clk,rst,matrix_A[868],matrix_B[68],mul_res1[868]);
multi_7x28 multi_7x28_mod_869(clk,rst,matrix_A[869],matrix_B[69],mul_res1[869]);
multi_7x28 multi_7x28_mod_870(clk,rst,matrix_A[870],matrix_B[70],mul_res1[870]);
multi_7x28 multi_7x28_mod_871(clk,rst,matrix_A[871],matrix_B[71],mul_res1[871]);
multi_7x28 multi_7x28_mod_872(clk,rst,matrix_A[872],matrix_B[72],mul_res1[872]);
multi_7x28 multi_7x28_mod_873(clk,rst,matrix_A[873],matrix_B[73],mul_res1[873]);
multi_7x28 multi_7x28_mod_874(clk,rst,matrix_A[874],matrix_B[74],mul_res1[874]);
multi_7x28 multi_7x28_mod_875(clk,rst,matrix_A[875],matrix_B[75],mul_res1[875]);
multi_7x28 multi_7x28_mod_876(clk,rst,matrix_A[876],matrix_B[76],mul_res1[876]);
multi_7x28 multi_7x28_mod_877(clk,rst,matrix_A[877],matrix_B[77],mul_res1[877]);
multi_7x28 multi_7x28_mod_878(clk,rst,matrix_A[878],matrix_B[78],mul_res1[878]);
multi_7x28 multi_7x28_mod_879(clk,rst,matrix_A[879],matrix_B[79],mul_res1[879]);
multi_7x28 multi_7x28_mod_880(clk,rst,matrix_A[880],matrix_B[80],mul_res1[880]);
multi_7x28 multi_7x28_mod_881(clk,rst,matrix_A[881],matrix_B[81],mul_res1[881]);
multi_7x28 multi_7x28_mod_882(clk,rst,matrix_A[882],matrix_B[82],mul_res1[882]);
multi_7x28 multi_7x28_mod_883(clk,rst,matrix_A[883],matrix_B[83],mul_res1[883]);
multi_7x28 multi_7x28_mod_884(clk,rst,matrix_A[884],matrix_B[84],mul_res1[884]);
multi_7x28 multi_7x28_mod_885(clk,rst,matrix_A[885],matrix_B[85],mul_res1[885]);
multi_7x28 multi_7x28_mod_886(clk,rst,matrix_A[886],matrix_B[86],mul_res1[886]);
multi_7x28 multi_7x28_mod_887(clk,rst,matrix_A[887],matrix_B[87],mul_res1[887]);
multi_7x28 multi_7x28_mod_888(clk,rst,matrix_A[888],matrix_B[88],mul_res1[888]);
multi_7x28 multi_7x28_mod_889(clk,rst,matrix_A[889],matrix_B[89],mul_res1[889]);
multi_7x28 multi_7x28_mod_890(clk,rst,matrix_A[890],matrix_B[90],mul_res1[890]);
multi_7x28 multi_7x28_mod_891(clk,rst,matrix_A[891],matrix_B[91],mul_res1[891]);
multi_7x28 multi_7x28_mod_892(clk,rst,matrix_A[892],matrix_B[92],mul_res1[892]);
multi_7x28 multi_7x28_mod_893(clk,rst,matrix_A[893],matrix_B[93],mul_res1[893]);
multi_7x28 multi_7x28_mod_894(clk,rst,matrix_A[894],matrix_B[94],mul_res1[894]);
multi_7x28 multi_7x28_mod_895(clk,rst,matrix_A[895],matrix_B[95],mul_res1[895]);
multi_7x28 multi_7x28_mod_896(clk,rst,matrix_A[896],matrix_B[96],mul_res1[896]);
multi_7x28 multi_7x28_mod_897(clk,rst,matrix_A[897],matrix_B[97],mul_res1[897]);
multi_7x28 multi_7x28_mod_898(clk,rst,matrix_A[898],matrix_B[98],mul_res1[898]);
multi_7x28 multi_7x28_mod_899(clk,rst,matrix_A[899],matrix_B[99],mul_res1[899]);
multi_7x28 multi_7x28_mod_900(clk,rst,matrix_A[900],matrix_B[100],mul_res1[900]);
multi_7x28 multi_7x28_mod_901(clk,rst,matrix_A[901],matrix_B[101],mul_res1[901]);
multi_7x28 multi_7x28_mod_902(clk,rst,matrix_A[902],matrix_B[102],mul_res1[902]);
multi_7x28 multi_7x28_mod_903(clk,rst,matrix_A[903],matrix_B[103],mul_res1[903]);
multi_7x28 multi_7x28_mod_904(clk,rst,matrix_A[904],matrix_B[104],mul_res1[904]);
multi_7x28 multi_7x28_mod_905(clk,rst,matrix_A[905],matrix_B[105],mul_res1[905]);
multi_7x28 multi_7x28_mod_906(clk,rst,matrix_A[906],matrix_B[106],mul_res1[906]);
multi_7x28 multi_7x28_mod_907(clk,rst,matrix_A[907],matrix_B[107],mul_res1[907]);
multi_7x28 multi_7x28_mod_908(clk,rst,matrix_A[908],matrix_B[108],mul_res1[908]);
multi_7x28 multi_7x28_mod_909(clk,rst,matrix_A[909],matrix_B[109],mul_res1[909]);
multi_7x28 multi_7x28_mod_910(clk,rst,matrix_A[910],matrix_B[110],mul_res1[910]);
multi_7x28 multi_7x28_mod_911(clk,rst,matrix_A[911],matrix_B[111],mul_res1[911]);
multi_7x28 multi_7x28_mod_912(clk,rst,matrix_A[912],matrix_B[112],mul_res1[912]);
multi_7x28 multi_7x28_mod_913(clk,rst,matrix_A[913],matrix_B[113],mul_res1[913]);
multi_7x28 multi_7x28_mod_914(clk,rst,matrix_A[914],matrix_B[114],mul_res1[914]);
multi_7x28 multi_7x28_mod_915(clk,rst,matrix_A[915],matrix_B[115],mul_res1[915]);
multi_7x28 multi_7x28_mod_916(clk,rst,matrix_A[916],matrix_B[116],mul_res1[916]);
multi_7x28 multi_7x28_mod_917(clk,rst,matrix_A[917],matrix_B[117],mul_res1[917]);
multi_7x28 multi_7x28_mod_918(clk,rst,matrix_A[918],matrix_B[118],mul_res1[918]);
multi_7x28 multi_7x28_mod_919(clk,rst,matrix_A[919],matrix_B[119],mul_res1[919]);
multi_7x28 multi_7x28_mod_920(clk,rst,matrix_A[920],matrix_B[120],mul_res1[920]);
multi_7x28 multi_7x28_mod_921(clk,rst,matrix_A[921],matrix_B[121],mul_res1[921]);
multi_7x28 multi_7x28_mod_922(clk,rst,matrix_A[922],matrix_B[122],mul_res1[922]);
multi_7x28 multi_7x28_mod_923(clk,rst,matrix_A[923],matrix_B[123],mul_res1[923]);
multi_7x28 multi_7x28_mod_924(clk,rst,matrix_A[924],matrix_B[124],mul_res1[924]);
multi_7x28 multi_7x28_mod_925(clk,rst,matrix_A[925],matrix_B[125],mul_res1[925]);
multi_7x28 multi_7x28_mod_926(clk,rst,matrix_A[926],matrix_B[126],mul_res1[926]);
multi_7x28 multi_7x28_mod_927(clk,rst,matrix_A[927],matrix_B[127],mul_res1[927]);
multi_7x28 multi_7x28_mod_928(clk,rst,matrix_A[928],matrix_B[128],mul_res1[928]);
multi_7x28 multi_7x28_mod_929(clk,rst,matrix_A[929],matrix_B[129],mul_res1[929]);
multi_7x28 multi_7x28_mod_930(clk,rst,matrix_A[930],matrix_B[130],mul_res1[930]);
multi_7x28 multi_7x28_mod_931(clk,rst,matrix_A[931],matrix_B[131],mul_res1[931]);
multi_7x28 multi_7x28_mod_932(clk,rst,matrix_A[932],matrix_B[132],mul_res1[932]);
multi_7x28 multi_7x28_mod_933(clk,rst,matrix_A[933],matrix_B[133],mul_res1[933]);
multi_7x28 multi_7x28_mod_934(clk,rst,matrix_A[934],matrix_B[134],mul_res1[934]);
multi_7x28 multi_7x28_mod_935(clk,rst,matrix_A[935],matrix_B[135],mul_res1[935]);
multi_7x28 multi_7x28_mod_936(clk,rst,matrix_A[936],matrix_B[136],mul_res1[936]);
multi_7x28 multi_7x28_mod_937(clk,rst,matrix_A[937],matrix_B[137],mul_res1[937]);
multi_7x28 multi_7x28_mod_938(clk,rst,matrix_A[938],matrix_B[138],mul_res1[938]);
multi_7x28 multi_7x28_mod_939(clk,rst,matrix_A[939],matrix_B[139],mul_res1[939]);
multi_7x28 multi_7x28_mod_940(clk,rst,matrix_A[940],matrix_B[140],mul_res1[940]);
multi_7x28 multi_7x28_mod_941(clk,rst,matrix_A[941],matrix_B[141],mul_res1[941]);
multi_7x28 multi_7x28_mod_942(clk,rst,matrix_A[942],matrix_B[142],mul_res1[942]);
multi_7x28 multi_7x28_mod_943(clk,rst,matrix_A[943],matrix_B[143],mul_res1[943]);
multi_7x28 multi_7x28_mod_944(clk,rst,matrix_A[944],matrix_B[144],mul_res1[944]);
multi_7x28 multi_7x28_mod_945(clk,rst,matrix_A[945],matrix_B[145],mul_res1[945]);
multi_7x28 multi_7x28_mod_946(clk,rst,matrix_A[946],matrix_B[146],mul_res1[946]);
multi_7x28 multi_7x28_mod_947(clk,rst,matrix_A[947],matrix_B[147],mul_res1[947]);
multi_7x28 multi_7x28_mod_948(clk,rst,matrix_A[948],matrix_B[148],mul_res1[948]);
multi_7x28 multi_7x28_mod_949(clk,rst,matrix_A[949],matrix_B[149],mul_res1[949]);
multi_7x28 multi_7x28_mod_950(clk,rst,matrix_A[950],matrix_B[150],mul_res1[950]);
multi_7x28 multi_7x28_mod_951(clk,rst,matrix_A[951],matrix_B[151],mul_res1[951]);
multi_7x28 multi_7x28_mod_952(clk,rst,matrix_A[952],matrix_B[152],mul_res1[952]);
multi_7x28 multi_7x28_mod_953(clk,rst,matrix_A[953],matrix_B[153],mul_res1[953]);
multi_7x28 multi_7x28_mod_954(clk,rst,matrix_A[954],matrix_B[154],mul_res1[954]);
multi_7x28 multi_7x28_mod_955(clk,rst,matrix_A[955],matrix_B[155],mul_res1[955]);
multi_7x28 multi_7x28_mod_956(clk,rst,matrix_A[956],matrix_B[156],mul_res1[956]);
multi_7x28 multi_7x28_mod_957(clk,rst,matrix_A[957],matrix_B[157],mul_res1[957]);
multi_7x28 multi_7x28_mod_958(clk,rst,matrix_A[958],matrix_B[158],mul_res1[958]);
multi_7x28 multi_7x28_mod_959(clk,rst,matrix_A[959],matrix_B[159],mul_res1[959]);
multi_7x28 multi_7x28_mod_960(clk,rst,matrix_A[960],matrix_B[160],mul_res1[960]);
multi_7x28 multi_7x28_mod_961(clk,rst,matrix_A[961],matrix_B[161],mul_res1[961]);
multi_7x28 multi_7x28_mod_962(clk,rst,matrix_A[962],matrix_B[162],mul_res1[962]);
multi_7x28 multi_7x28_mod_963(clk,rst,matrix_A[963],matrix_B[163],mul_res1[963]);
multi_7x28 multi_7x28_mod_964(clk,rst,matrix_A[964],matrix_B[164],mul_res1[964]);
multi_7x28 multi_7x28_mod_965(clk,rst,matrix_A[965],matrix_B[165],mul_res1[965]);
multi_7x28 multi_7x28_mod_966(clk,rst,matrix_A[966],matrix_B[166],mul_res1[966]);
multi_7x28 multi_7x28_mod_967(clk,rst,matrix_A[967],matrix_B[167],mul_res1[967]);
multi_7x28 multi_7x28_mod_968(clk,rst,matrix_A[968],matrix_B[168],mul_res1[968]);
multi_7x28 multi_7x28_mod_969(clk,rst,matrix_A[969],matrix_B[169],mul_res1[969]);
multi_7x28 multi_7x28_mod_970(clk,rst,matrix_A[970],matrix_B[170],mul_res1[970]);
multi_7x28 multi_7x28_mod_971(clk,rst,matrix_A[971],matrix_B[171],mul_res1[971]);
multi_7x28 multi_7x28_mod_972(clk,rst,matrix_A[972],matrix_B[172],mul_res1[972]);
multi_7x28 multi_7x28_mod_973(clk,rst,matrix_A[973],matrix_B[173],mul_res1[973]);
multi_7x28 multi_7x28_mod_974(clk,rst,matrix_A[974],matrix_B[174],mul_res1[974]);
multi_7x28 multi_7x28_mod_975(clk,rst,matrix_A[975],matrix_B[175],mul_res1[975]);
multi_7x28 multi_7x28_mod_976(clk,rst,matrix_A[976],matrix_B[176],mul_res1[976]);
multi_7x28 multi_7x28_mod_977(clk,rst,matrix_A[977],matrix_B[177],mul_res1[977]);
multi_7x28 multi_7x28_mod_978(clk,rst,matrix_A[978],matrix_B[178],mul_res1[978]);
multi_7x28 multi_7x28_mod_979(clk,rst,matrix_A[979],matrix_B[179],mul_res1[979]);
multi_7x28 multi_7x28_mod_980(clk,rst,matrix_A[980],matrix_B[180],mul_res1[980]);
multi_7x28 multi_7x28_mod_981(clk,rst,matrix_A[981],matrix_B[181],mul_res1[981]);
multi_7x28 multi_7x28_mod_982(clk,rst,matrix_A[982],matrix_B[182],mul_res1[982]);
multi_7x28 multi_7x28_mod_983(clk,rst,matrix_A[983],matrix_B[183],mul_res1[983]);
multi_7x28 multi_7x28_mod_984(clk,rst,matrix_A[984],matrix_B[184],mul_res1[984]);
multi_7x28 multi_7x28_mod_985(clk,rst,matrix_A[985],matrix_B[185],mul_res1[985]);
multi_7x28 multi_7x28_mod_986(clk,rst,matrix_A[986],matrix_B[186],mul_res1[986]);
multi_7x28 multi_7x28_mod_987(clk,rst,matrix_A[987],matrix_B[187],mul_res1[987]);
multi_7x28 multi_7x28_mod_988(clk,rst,matrix_A[988],matrix_B[188],mul_res1[988]);
multi_7x28 multi_7x28_mod_989(clk,rst,matrix_A[989],matrix_B[189],mul_res1[989]);
multi_7x28 multi_7x28_mod_990(clk,rst,matrix_A[990],matrix_B[190],mul_res1[990]);
multi_7x28 multi_7x28_mod_991(clk,rst,matrix_A[991],matrix_B[191],mul_res1[991]);
multi_7x28 multi_7x28_mod_992(clk,rst,matrix_A[992],matrix_B[192],mul_res1[992]);
multi_7x28 multi_7x28_mod_993(clk,rst,matrix_A[993],matrix_B[193],mul_res1[993]);
multi_7x28 multi_7x28_mod_994(clk,rst,matrix_A[994],matrix_B[194],mul_res1[994]);
multi_7x28 multi_7x28_mod_995(clk,rst,matrix_A[995],matrix_B[195],mul_res1[995]);
multi_7x28 multi_7x28_mod_996(clk,rst,matrix_A[996],matrix_B[196],mul_res1[996]);
multi_7x28 multi_7x28_mod_997(clk,rst,matrix_A[997],matrix_B[197],mul_res1[997]);
multi_7x28 multi_7x28_mod_998(clk,rst,matrix_A[998],matrix_B[198],mul_res1[998]);
multi_7x28 multi_7x28_mod_999(clk,rst,matrix_A[999],matrix_B[199],mul_res1[999]);
multi_7x28 multi_7x28_mod_1000(clk,rst,matrix_A[1000],matrix_B[0],mul_res1[1000]);
multi_7x28 multi_7x28_mod_1001(clk,rst,matrix_A[1001],matrix_B[1],mul_res1[1001]);
multi_7x28 multi_7x28_mod_1002(clk,rst,matrix_A[1002],matrix_B[2],mul_res1[1002]);
multi_7x28 multi_7x28_mod_1003(clk,rst,matrix_A[1003],matrix_B[3],mul_res1[1003]);
multi_7x28 multi_7x28_mod_1004(clk,rst,matrix_A[1004],matrix_B[4],mul_res1[1004]);
multi_7x28 multi_7x28_mod_1005(clk,rst,matrix_A[1005],matrix_B[5],mul_res1[1005]);
multi_7x28 multi_7x28_mod_1006(clk,rst,matrix_A[1006],matrix_B[6],mul_res1[1006]);
multi_7x28 multi_7x28_mod_1007(clk,rst,matrix_A[1007],matrix_B[7],mul_res1[1007]);
multi_7x28 multi_7x28_mod_1008(clk,rst,matrix_A[1008],matrix_B[8],mul_res1[1008]);
multi_7x28 multi_7x28_mod_1009(clk,rst,matrix_A[1009],matrix_B[9],mul_res1[1009]);
multi_7x28 multi_7x28_mod_1010(clk,rst,matrix_A[1010],matrix_B[10],mul_res1[1010]);
multi_7x28 multi_7x28_mod_1011(clk,rst,matrix_A[1011],matrix_B[11],mul_res1[1011]);
multi_7x28 multi_7x28_mod_1012(clk,rst,matrix_A[1012],matrix_B[12],mul_res1[1012]);
multi_7x28 multi_7x28_mod_1013(clk,rst,matrix_A[1013],matrix_B[13],mul_res1[1013]);
multi_7x28 multi_7x28_mod_1014(clk,rst,matrix_A[1014],matrix_B[14],mul_res1[1014]);
multi_7x28 multi_7x28_mod_1015(clk,rst,matrix_A[1015],matrix_B[15],mul_res1[1015]);
multi_7x28 multi_7x28_mod_1016(clk,rst,matrix_A[1016],matrix_B[16],mul_res1[1016]);
multi_7x28 multi_7x28_mod_1017(clk,rst,matrix_A[1017],matrix_B[17],mul_res1[1017]);
multi_7x28 multi_7x28_mod_1018(clk,rst,matrix_A[1018],matrix_B[18],mul_res1[1018]);
multi_7x28 multi_7x28_mod_1019(clk,rst,matrix_A[1019],matrix_B[19],mul_res1[1019]);
multi_7x28 multi_7x28_mod_1020(clk,rst,matrix_A[1020],matrix_B[20],mul_res1[1020]);
multi_7x28 multi_7x28_mod_1021(clk,rst,matrix_A[1021],matrix_B[21],mul_res1[1021]);
multi_7x28 multi_7x28_mod_1022(clk,rst,matrix_A[1022],matrix_B[22],mul_res1[1022]);
multi_7x28 multi_7x28_mod_1023(clk,rst,matrix_A[1023],matrix_B[23],mul_res1[1023]);
multi_7x28 multi_7x28_mod_1024(clk,rst,matrix_A[1024],matrix_B[24],mul_res1[1024]);
multi_7x28 multi_7x28_mod_1025(clk,rst,matrix_A[1025],matrix_B[25],mul_res1[1025]);
multi_7x28 multi_7x28_mod_1026(clk,rst,matrix_A[1026],matrix_B[26],mul_res1[1026]);
multi_7x28 multi_7x28_mod_1027(clk,rst,matrix_A[1027],matrix_B[27],mul_res1[1027]);
multi_7x28 multi_7x28_mod_1028(clk,rst,matrix_A[1028],matrix_B[28],mul_res1[1028]);
multi_7x28 multi_7x28_mod_1029(clk,rst,matrix_A[1029],matrix_B[29],mul_res1[1029]);
multi_7x28 multi_7x28_mod_1030(clk,rst,matrix_A[1030],matrix_B[30],mul_res1[1030]);
multi_7x28 multi_7x28_mod_1031(clk,rst,matrix_A[1031],matrix_B[31],mul_res1[1031]);
multi_7x28 multi_7x28_mod_1032(clk,rst,matrix_A[1032],matrix_B[32],mul_res1[1032]);
multi_7x28 multi_7x28_mod_1033(clk,rst,matrix_A[1033],matrix_B[33],mul_res1[1033]);
multi_7x28 multi_7x28_mod_1034(clk,rst,matrix_A[1034],matrix_B[34],mul_res1[1034]);
multi_7x28 multi_7x28_mod_1035(clk,rst,matrix_A[1035],matrix_B[35],mul_res1[1035]);
multi_7x28 multi_7x28_mod_1036(clk,rst,matrix_A[1036],matrix_B[36],mul_res1[1036]);
multi_7x28 multi_7x28_mod_1037(clk,rst,matrix_A[1037],matrix_B[37],mul_res1[1037]);
multi_7x28 multi_7x28_mod_1038(clk,rst,matrix_A[1038],matrix_B[38],mul_res1[1038]);
multi_7x28 multi_7x28_mod_1039(clk,rst,matrix_A[1039],matrix_B[39],mul_res1[1039]);
multi_7x28 multi_7x28_mod_1040(clk,rst,matrix_A[1040],matrix_B[40],mul_res1[1040]);
multi_7x28 multi_7x28_mod_1041(clk,rst,matrix_A[1041],matrix_B[41],mul_res1[1041]);
multi_7x28 multi_7x28_mod_1042(clk,rst,matrix_A[1042],matrix_B[42],mul_res1[1042]);
multi_7x28 multi_7x28_mod_1043(clk,rst,matrix_A[1043],matrix_B[43],mul_res1[1043]);
multi_7x28 multi_7x28_mod_1044(clk,rst,matrix_A[1044],matrix_B[44],mul_res1[1044]);
multi_7x28 multi_7x28_mod_1045(clk,rst,matrix_A[1045],matrix_B[45],mul_res1[1045]);
multi_7x28 multi_7x28_mod_1046(clk,rst,matrix_A[1046],matrix_B[46],mul_res1[1046]);
multi_7x28 multi_7x28_mod_1047(clk,rst,matrix_A[1047],matrix_B[47],mul_res1[1047]);
multi_7x28 multi_7x28_mod_1048(clk,rst,matrix_A[1048],matrix_B[48],mul_res1[1048]);
multi_7x28 multi_7x28_mod_1049(clk,rst,matrix_A[1049],matrix_B[49],mul_res1[1049]);
multi_7x28 multi_7x28_mod_1050(clk,rst,matrix_A[1050],matrix_B[50],mul_res1[1050]);
multi_7x28 multi_7x28_mod_1051(clk,rst,matrix_A[1051],matrix_B[51],mul_res1[1051]);
multi_7x28 multi_7x28_mod_1052(clk,rst,matrix_A[1052],matrix_B[52],mul_res1[1052]);
multi_7x28 multi_7x28_mod_1053(clk,rst,matrix_A[1053],matrix_B[53],mul_res1[1053]);
multi_7x28 multi_7x28_mod_1054(clk,rst,matrix_A[1054],matrix_B[54],mul_res1[1054]);
multi_7x28 multi_7x28_mod_1055(clk,rst,matrix_A[1055],matrix_B[55],mul_res1[1055]);
multi_7x28 multi_7x28_mod_1056(clk,rst,matrix_A[1056],matrix_B[56],mul_res1[1056]);
multi_7x28 multi_7x28_mod_1057(clk,rst,matrix_A[1057],matrix_B[57],mul_res1[1057]);
multi_7x28 multi_7x28_mod_1058(clk,rst,matrix_A[1058],matrix_B[58],mul_res1[1058]);
multi_7x28 multi_7x28_mod_1059(clk,rst,matrix_A[1059],matrix_B[59],mul_res1[1059]);
multi_7x28 multi_7x28_mod_1060(clk,rst,matrix_A[1060],matrix_B[60],mul_res1[1060]);
multi_7x28 multi_7x28_mod_1061(clk,rst,matrix_A[1061],matrix_B[61],mul_res1[1061]);
multi_7x28 multi_7x28_mod_1062(clk,rst,matrix_A[1062],matrix_B[62],mul_res1[1062]);
multi_7x28 multi_7x28_mod_1063(clk,rst,matrix_A[1063],matrix_B[63],mul_res1[1063]);
multi_7x28 multi_7x28_mod_1064(clk,rst,matrix_A[1064],matrix_B[64],mul_res1[1064]);
multi_7x28 multi_7x28_mod_1065(clk,rst,matrix_A[1065],matrix_B[65],mul_res1[1065]);
multi_7x28 multi_7x28_mod_1066(clk,rst,matrix_A[1066],matrix_B[66],mul_res1[1066]);
multi_7x28 multi_7x28_mod_1067(clk,rst,matrix_A[1067],matrix_B[67],mul_res1[1067]);
multi_7x28 multi_7x28_mod_1068(clk,rst,matrix_A[1068],matrix_B[68],mul_res1[1068]);
multi_7x28 multi_7x28_mod_1069(clk,rst,matrix_A[1069],matrix_B[69],mul_res1[1069]);
multi_7x28 multi_7x28_mod_1070(clk,rst,matrix_A[1070],matrix_B[70],mul_res1[1070]);
multi_7x28 multi_7x28_mod_1071(clk,rst,matrix_A[1071],matrix_B[71],mul_res1[1071]);
multi_7x28 multi_7x28_mod_1072(clk,rst,matrix_A[1072],matrix_B[72],mul_res1[1072]);
multi_7x28 multi_7x28_mod_1073(clk,rst,matrix_A[1073],matrix_B[73],mul_res1[1073]);
multi_7x28 multi_7x28_mod_1074(clk,rst,matrix_A[1074],matrix_B[74],mul_res1[1074]);
multi_7x28 multi_7x28_mod_1075(clk,rst,matrix_A[1075],matrix_B[75],mul_res1[1075]);
multi_7x28 multi_7x28_mod_1076(clk,rst,matrix_A[1076],matrix_B[76],mul_res1[1076]);
multi_7x28 multi_7x28_mod_1077(clk,rst,matrix_A[1077],matrix_B[77],mul_res1[1077]);
multi_7x28 multi_7x28_mod_1078(clk,rst,matrix_A[1078],matrix_B[78],mul_res1[1078]);
multi_7x28 multi_7x28_mod_1079(clk,rst,matrix_A[1079],matrix_B[79],mul_res1[1079]);
multi_7x28 multi_7x28_mod_1080(clk,rst,matrix_A[1080],matrix_B[80],mul_res1[1080]);
multi_7x28 multi_7x28_mod_1081(clk,rst,matrix_A[1081],matrix_B[81],mul_res1[1081]);
multi_7x28 multi_7x28_mod_1082(clk,rst,matrix_A[1082],matrix_B[82],mul_res1[1082]);
multi_7x28 multi_7x28_mod_1083(clk,rst,matrix_A[1083],matrix_B[83],mul_res1[1083]);
multi_7x28 multi_7x28_mod_1084(clk,rst,matrix_A[1084],matrix_B[84],mul_res1[1084]);
multi_7x28 multi_7x28_mod_1085(clk,rst,matrix_A[1085],matrix_B[85],mul_res1[1085]);
multi_7x28 multi_7x28_mod_1086(clk,rst,matrix_A[1086],matrix_B[86],mul_res1[1086]);
multi_7x28 multi_7x28_mod_1087(clk,rst,matrix_A[1087],matrix_B[87],mul_res1[1087]);
multi_7x28 multi_7x28_mod_1088(clk,rst,matrix_A[1088],matrix_B[88],mul_res1[1088]);
multi_7x28 multi_7x28_mod_1089(clk,rst,matrix_A[1089],matrix_B[89],mul_res1[1089]);
multi_7x28 multi_7x28_mod_1090(clk,rst,matrix_A[1090],matrix_B[90],mul_res1[1090]);
multi_7x28 multi_7x28_mod_1091(clk,rst,matrix_A[1091],matrix_B[91],mul_res1[1091]);
multi_7x28 multi_7x28_mod_1092(clk,rst,matrix_A[1092],matrix_B[92],mul_res1[1092]);
multi_7x28 multi_7x28_mod_1093(clk,rst,matrix_A[1093],matrix_B[93],mul_res1[1093]);
multi_7x28 multi_7x28_mod_1094(clk,rst,matrix_A[1094],matrix_B[94],mul_res1[1094]);
multi_7x28 multi_7x28_mod_1095(clk,rst,matrix_A[1095],matrix_B[95],mul_res1[1095]);
multi_7x28 multi_7x28_mod_1096(clk,rst,matrix_A[1096],matrix_B[96],mul_res1[1096]);
multi_7x28 multi_7x28_mod_1097(clk,rst,matrix_A[1097],matrix_B[97],mul_res1[1097]);
multi_7x28 multi_7x28_mod_1098(clk,rst,matrix_A[1098],matrix_B[98],mul_res1[1098]);
multi_7x28 multi_7x28_mod_1099(clk,rst,matrix_A[1099],matrix_B[99],mul_res1[1099]);
multi_7x28 multi_7x28_mod_1100(clk,rst,matrix_A[1100],matrix_B[100],mul_res1[1100]);
multi_7x28 multi_7x28_mod_1101(clk,rst,matrix_A[1101],matrix_B[101],mul_res1[1101]);
multi_7x28 multi_7x28_mod_1102(clk,rst,matrix_A[1102],matrix_B[102],mul_res1[1102]);
multi_7x28 multi_7x28_mod_1103(clk,rst,matrix_A[1103],matrix_B[103],mul_res1[1103]);
multi_7x28 multi_7x28_mod_1104(clk,rst,matrix_A[1104],matrix_B[104],mul_res1[1104]);
multi_7x28 multi_7x28_mod_1105(clk,rst,matrix_A[1105],matrix_B[105],mul_res1[1105]);
multi_7x28 multi_7x28_mod_1106(clk,rst,matrix_A[1106],matrix_B[106],mul_res1[1106]);
multi_7x28 multi_7x28_mod_1107(clk,rst,matrix_A[1107],matrix_B[107],mul_res1[1107]);
multi_7x28 multi_7x28_mod_1108(clk,rst,matrix_A[1108],matrix_B[108],mul_res1[1108]);
multi_7x28 multi_7x28_mod_1109(clk,rst,matrix_A[1109],matrix_B[109],mul_res1[1109]);
multi_7x28 multi_7x28_mod_1110(clk,rst,matrix_A[1110],matrix_B[110],mul_res1[1110]);
multi_7x28 multi_7x28_mod_1111(clk,rst,matrix_A[1111],matrix_B[111],mul_res1[1111]);
multi_7x28 multi_7x28_mod_1112(clk,rst,matrix_A[1112],matrix_B[112],mul_res1[1112]);
multi_7x28 multi_7x28_mod_1113(clk,rst,matrix_A[1113],matrix_B[113],mul_res1[1113]);
multi_7x28 multi_7x28_mod_1114(clk,rst,matrix_A[1114],matrix_B[114],mul_res1[1114]);
multi_7x28 multi_7x28_mod_1115(clk,rst,matrix_A[1115],matrix_B[115],mul_res1[1115]);
multi_7x28 multi_7x28_mod_1116(clk,rst,matrix_A[1116],matrix_B[116],mul_res1[1116]);
multi_7x28 multi_7x28_mod_1117(clk,rst,matrix_A[1117],matrix_B[117],mul_res1[1117]);
multi_7x28 multi_7x28_mod_1118(clk,rst,matrix_A[1118],matrix_B[118],mul_res1[1118]);
multi_7x28 multi_7x28_mod_1119(clk,rst,matrix_A[1119],matrix_B[119],mul_res1[1119]);
multi_7x28 multi_7x28_mod_1120(clk,rst,matrix_A[1120],matrix_B[120],mul_res1[1120]);
multi_7x28 multi_7x28_mod_1121(clk,rst,matrix_A[1121],matrix_B[121],mul_res1[1121]);
multi_7x28 multi_7x28_mod_1122(clk,rst,matrix_A[1122],matrix_B[122],mul_res1[1122]);
multi_7x28 multi_7x28_mod_1123(clk,rst,matrix_A[1123],matrix_B[123],mul_res1[1123]);
multi_7x28 multi_7x28_mod_1124(clk,rst,matrix_A[1124],matrix_B[124],mul_res1[1124]);
multi_7x28 multi_7x28_mod_1125(clk,rst,matrix_A[1125],matrix_B[125],mul_res1[1125]);
multi_7x28 multi_7x28_mod_1126(clk,rst,matrix_A[1126],matrix_B[126],mul_res1[1126]);
multi_7x28 multi_7x28_mod_1127(clk,rst,matrix_A[1127],matrix_B[127],mul_res1[1127]);
multi_7x28 multi_7x28_mod_1128(clk,rst,matrix_A[1128],matrix_B[128],mul_res1[1128]);
multi_7x28 multi_7x28_mod_1129(clk,rst,matrix_A[1129],matrix_B[129],mul_res1[1129]);
multi_7x28 multi_7x28_mod_1130(clk,rst,matrix_A[1130],matrix_B[130],mul_res1[1130]);
multi_7x28 multi_7x28_mod_1131(clk,rst,matrix_A[1131],matrix_B[131],mul_res1[1131]);
multi_7x28 multi_7x28_mod_1132(clk,rst,matrix_A[1132],matrix_B[132],mul_res1[1132]);
multi_7x28 multi_7x28_mod_1133(clk,rst,matrix_A[1133],matrix_B[133],mul_res1[1133]);
multi_7x28 multi_7x28_mod_1134(clk,rst,matrix_A[1134],matrix_B[134],mul_res1[1134]);
multi_7x28 multi_7x28_mod_1135(clk,rst,matrix_A[1135],matrix_B[135],mul_res1[1135]);
multi_7x28 multi_7x28_mod_1136(clk,rst,matrix_A[1136],matrix_B[136],mul_res1[1136]);
multi_7x28 multi_7x28_mod_1137(clk,rst,matrix_A[1137],matrix_B[137],mul_res1[1137]);
multi_7x28 multi_7x28_mod_1138(clk,rst,matrix_A[1138],matrix_B[138],mul_res1[1138]);
multi_7x28 multi_7x28_mod_1139(clk,rst,matrix_A[1139],matrix_B[139],mul_res1[1139]);
multi_7x28 multi_7x28_mod_1140(clk,rst,matrix_A[1140],matrix_B[140],mul_res1[1140]);
multi_7x28 multi_7x28_mod_1141(clk,rst,matrix_A[1141],matrix_B[141],mul_res1[1141]);
multi_7x28 multi_7x28_mod_1142(clk,rst,matrix_A[1142],matrix_B[142],mul_res1[1142]);
multi_7x28 multi_7x28_mod_1143(clk,rst,matrix_A[1143],matrix_B[143],mul_res1[1143]);
multi_7x28 multi_7x28_mod_1144(clk,rst,matrix_A[1144],matrix_B[144],mul_res1[1144]);
multi_7x28 multi_7x28_mod_1145(clk,rst,matrix_A[1145],matrix_B[145],mul_res1[1145]);
multi_7x28 multi_7x28_mod_1146(clk,rst,matrix_A[1146],matrix_B[146],mul_res1[1146]);
multi_7x28 multi_7x28_mod_1147(clk,rst,matrix_A[1147],matrix_B[147],mul_res1[1147]);
multi_7x28 multi_7x28_mod_1148(clk,rst,matrix_A[1148],matrix_B[148],mul_res1[1148]);
multi_7x28 multi_7x28_mod_1149(clk,rst,matrix_A[1149],matrix_B[149],mul_res1[1149]);
multi_7x28 multi_7x28_mod_1150(clk,rst,matrix_A[1150],matrix_B[150],mul_res1[1150]);
multi_7x28 multi_7x28_mod_1151(clk,rst,matrix_A[1151],matrix_B[151],mul_res1[1151]);
multi_7x28 multi_7x28_mod_1152(clk,rst,matrix_A[1152],matrix_B[152],mul_res1[1152]);
multi_7x28 multi_7x28_mod_1153(clk,rst,matrix_A[1153],matrix_B[153],mul_res1[1153]);
multi_7x28 multi_7x28_mod_1154(clk,rst,matrix_A[1154],matrix_B[154],mul_res1[1154]);
multi_7x28 multi_7x28_mod_1155(clk,rst,matrix_A[1155],matrix_B[155],mul_res1[1155]);
multi_7x28 multi_7x28_mod_1156(clk,rst,matrix_A[1156],matrix_B[156],mul_res1[1156]);
multi_7x28 multi_7x28_mod_1157(clk,rst,matrix_A[1157],matrix_B[157],mul_res1[1157]);
multi_7x28 multi_7x28_mod_1158(clk,rst,matrix_A[1158],matrix_B[158],mul_res1[1158]);
multi_7x28 multi_7x28_mod_1159(clk,rst,matrix_A[1159],matrix_B[159],mul_res1[1159]);
multi_7x28 multi_7x28_mod_1160(clk,rst,matrix_A[1160],matrix_B[160],mul_res1[1160]);
multi_7x28 multi_7x28_mod_1161(clk,rst,matrix_A[1161],matrix_B[161],mul_res1[1161]);
multi_7x28 multi_7x28_mod_1162(clk,rst,matrix_A[1162],matrix_B[162],mul_res1[1162]);
multi_7x28 multi_7x28_mod_1163(clk,rst,matrix_A[1163],matrix_B[163],mul_res1[1163]);
multi_7x28 multi_7x28_mod_1164(clk,rst,matrix_A[1164],matrix_B[164],mul_res1[1164]);
multi_7x28 multi_7x28_mod_1165(clk,rst,matrix_A[1165],matrix_B[165],mul_res1[1165]);
multi_7x28 multi_7x28_mod_1166(clk,rst,matrix_A[1166],matrix_B[166],mul_res1[1166]);
multi_7x28 multi_7x28_mod_1167(clk,rst,matrix_A[1167],matrix_B[167],mul_res1[1167]);
multi_7x28 multi_7x28_mod_1168(clk,rst,matrix_A[1168],matrix_B[168],mul_res1[1168]);
multi_7x28 multi_7x28_mod_1169(clk,rst,matrix_A[1169],matrix_B[169],mul_res1[1169]);
multi_7x28 multi_7x28_mod_1170(clk,rst,matrix_A[1170],matrix_B[170],mul_res1[1170]);
multi_7x28 multi_7x28_mod_1171(clk,rst,matrix_A[1171],matrix_B[171],mul_res1[1171]);
multi_7x28 multi_7x28_mod_1172(clk,rst,matrix_A[1172],matrix_B[172],mul_res1[1172]);
multi_7x28 multi_7x28_mod_1173(clk,rst,matrix_A[1173],matrix_B[173],mul_res1[1173]);
multi_7x28 multi_7x28_mod_1174(clk,rst,matrix_A[1174],matrix_B[174],mul_res1[1174]);
multi_7x28 multi_7x28_mod_1175(clk,rst,matrix_A[1175],matrix_B[175],mul_res1[1175]);
multi_7x28 multi_7x28_mod_1176(clk,rst,matrix_A[1176],matrix_B[176],mul_res1[1176]);
multi_7x28 multi_7x28_mod_1177(clk,rst,matrix_A[1177],matrix_B[177],mul_res1[1177]);
multi_7x28 multi_7x28_mod_1178(clk,rst,matrix_A[1178],matrix_B[178],mul_res1[1178]);
multi_7x28 multi_7x28_mod_1179(clk,rst,matrix_A[1179],matrix_B[179],mul_res1[1179]);
multi_7x28 multi_7x28_mod_1180(clk,rst,matrix_A[1180],matrix_B[180],mul_res1[1180]);
multi_7x28 multi_7x28_mod_1181(clk,rst,matrix_A[1181],matrix_B[181],mul_res1[1181]);
multi_7x28 multi_7x28_mod_1182(clk,rst,matrix_A[1182],matrix_B[182],mul_res1[1182]);
multi_7x28 multi_7x28_mod_1183(clk,rst,matrix_A[1183],matrix_B[183],mul_res1[1183]);
multi_7x28 multi_7x28_mod_1184(clk,rst,matrix_A[1184],matrix_B[184],mul_res1[1184]);
multi_7x28 multi_7x28_mod_1185(clk,rst,matrix_A[1185],matrix_B[185],mul_res1[1185]);
multi_7x28 multi_7x28_mod_1186(clk,rst,matrix_A[1186],matrix_B[186],mul_res1[1186]);
multi_7x28 multi_7x28_mod_1187(clk,rst,matrix_A[1187],matrix_B[187],mul_res1[1187]);
multi_7x28 multi_7x28_mod_1188(clk,rst,matrix_A[1188],matrix_B[188],mul_res1[1188]);
multi_7x28 multi_7x28_mod_1189(clk,rst,matrix_A[1189],matrix_B[189],mul_res1[1189]);
multi_7x28 multi_7x28_mod_1190(clk,rst,matrix_A[1190],matrix_B[190],mul_res1[1190]);
multi_7x28 multi_7x28_mod_1191(clk,rst,matrix_A[1191],matrix_B[191],mul_res1[1191]);
multi_7x28 multi_7x28_mod_1192(clk,rst,matrix_A[1192],matrix_B[192],mul_res1[1192]);
multi_7x28 multi_7x28_mod_1193(clk,rst,matrix_A[1193],matrix_B[193],mul_res1[1193]);
multi_7x28 multi_7x28_mod_1194(clk,rst,matrix_A[1194],matrix_B[194],mul_res1[1194]);
multi_7x28 multi_7x28_mod_1195(clk,rst,matrix_A[1195],matrix_B[195],mul_res1[1195]);
multi_7x28 multi_7x28_mod_1196(clk,rst,matrix_A[1196],matrix_B[196],mul_res1[1196]);
multi_7x28 multi_7x28_mod_1197(clk,rst,matrix_A[1197],matrix_B[197],mul_res1[1197]);
multi_7x28 multi_7x28_mod_1198(clk,rst,matrix_A[1198],matrix_B[198],mul_res1[1198]);
multi_7x28 multi_7x28_mod_1199(clk,rst,matrix_A[1199],matrix_B[199],mul_res1[1199]);
multi_7x28 multi_7x28_mod_1200(clk,rst,matrix_A[1200],matrix_B[0],mul_res1[1200]);
multi_7x28 multi_7x28_mod_1201(clk,rst,matrix_A[1201],matrix_B[1],mul_res1[1201]);
multi_7x28 multi_7x28_mod_1202(clk,rst,matrix_A[1202],matrix_B[2],mul_res1[1202]);
multi_7x28 multi_7x28_mod_1203(clk,rst,matrix_A[1203],matrix_B[3],mul_res1[1203]);
multi_7x28 multi_7x28_mod_1204(clk,rst,matrix_A[1204],matrix_B[4],mul_res1[1204]);
multi_7x28 multi_7x28_mod_1205(clk,rst,matrix_A[1205],matrix_B[5],mul_res1[1205]);
multi_7x28 multi_7x28_mod_1206(clk,rst,matrix_A[1206],matrix_B[6],mul_res1[1206]);
multi_7x28 multi_7x28_mod_1207(clk,rst,matrix_A[1207],matrix_B[7],mul_res1[1207]);
multi_7x28 multi_7x28_mod_1208(clk,rst,matrix_A[1208],matrix_B[8],mul_res1[1208]);
multi_7x28 multi_7x28_mod_1209(clk,rst,matrix_A[1209],matrix_B[9],mul_res1[1209]);
multi_7x28 multi_7x28_mod_1210(clk,rst,matrix_A[1210],matrix_B[10],mul_res1[1210]);
multi_7x28 multi_7x28_mod_1211(clk,rst,matrix_A[1211],matrix_B[11],mul_res1[1211]);
multi_7x28 multi_7x28_mod_1212(clk,rst,matrix_A[1212],matrix_B[12],mul_res1[1212]);
multi_7x28 multi_7x28_mod_1213(clk,rst,matrix_A[1213],matrix_B[13],mul_res1[1213]);
multi_7x28 multi_7x28_mod_1214(clk,rst,matrix_A[1214],matrix_B[14],mul_res1[1214]);
multi_7x28 multi_7x28_mod_1215(clk,rst,matrix_A[1215],matrix_B[15],mul_res1[1215]);
multi_7x28 multi_7x28_mod_1216(clk,rst,matrix_A[1216],matrix_B[16],mul_res1[1216]);
multi_7x28 multi_7x28_mod_1217(clk,rst,matrix_A[1217],matrix_B[17],mul_res1[1217]);
multi_7x28 multi_7x28_mod_1218(clk,rst,matrix_A[1218],matrix_B[18],mul_res1[1218]);
multi_7x28 multi_7x28_mod_1219(clk,rst,matrix_A[1219],matrix_B[19],mul_res1[1219]);
multi_7x28 multi_7x28_mod_1220(clk,rst,matrix_A[1220],matrix_B[20],mul_res1[1220]);
multi_7x28 multi_7x28_mod_1221(clk,rst,matrix_A[1221],matrix_B[21],mul_res1[1221]);
multi_7x28 multi_7x28_mod_1222(clk,rst,matrix_A[1222],matrix_B[22],mul_res1[1222]);
multi_7x28 multi_7x28_mod_1223(clk,rst,matrix_A[1223],matrix_B[23],mul_res1[1223]);
multi_7x28 multi_7x28_mod_1224(clk,rst,matrix_A[1224],matrix_B[24],mul_res1[1224]);
multi_7x28 multi_7x28_mod_1225(clk,rst,matrix_A[1225],matrix_B[25],mul_res1[1225]);
multi_7x28 multi_7x28_mod_1226(clk,rst,matrix_A[1226],matrix_B[26],mul_res1[1226]);
multi_7x28 multi_7x28_mod_1227(clk,rst,matrix_A[1227],matrix_B[27],mul_res1[1227]);
multi_7x28 multi_7x28_mod_1228(clk,rst,matrix_A[1228],matrix_B[28],mul_res1[1228]);
multi_7x28 multi_7x28_mod_1229(clk,rst,matrix_A[1229],matrix_B[29],mul_res1[1229]);
multi_7x28 multi_7x28_mod_1230(clk,rst,matrix_A[1230],matrix_B[30],mul_res1[1230]);
multi_7x28 multi_7x28_mod_1231(clk,rst,matrix_A[1231],matrix_B[31],mul_res1[1231]);
multi_7x28 multi_7x28_mod_1232(clk,rst,matrix_A[1232],matrix_B[32],mul_res1[1232]);
multi_7x28 multi_7x28_mod_1233(clk,rst,matrix_A[1233],matrix_B[33],mul_res1[1233]);
multi_7x28 multi_7x28_mod_1234(clk,rst,matrix_A[1234],matrix_B[34],mul_res1[1234]);
multi_7x28 multi_7x28_mod_1235(clk,rst,matrix_A[1235],matrix_B[35],mul_res1[1235]);
multi_7x28 multi_7x28_mod_1236(clk,rst,matrix_A[1236],matrix_B[36],mul_res1[1236]);
multi_7x28 multi_7x28_mod_1237(clk,rst,matrix_A[1237],matrix_B[37],mul_res1[1237]);
multi_7x28 multi_7x28_mod_1238(clk,rst,matrix_A[1238],matrix_B[38],mul_res1[1238]);
multi_7x28 multi_7x28_mod_1239(clk,rst,matrix_A[1239],matrix_B[39],mul_res1[1239]);
multi_7x28 multi_7x28_mod_1240(clk,rst,matrix_A[1240],matrix_B[40],mul_res1[1240]);
multi_7x28 multi_7x28_mod_1241(clk,rst,matrix_A[1241],matrix_B[41],mul_res1[1241]);
multi_7x28 multi_7x28_mod_1242(clk,rst,matrix_A[1242],matrix_B[42],mul_res1[1242]);
multi_7x28 multi_7x28_mod_1243(clk,rst,matrix_A[1243],matrix_B[43],mul_res1[1243]);
multi_7x28 multi_7x28_mod_1244(clk,rst,matrix_A[1244],matrix_B[44],mul_res1[1244]);
multi_7x28 multi_7x28_mod_1245(clk,rst,matrix_A[1245],matrix_B[45],mul_res1[1245]);
multi_7x28 multi_7x28_mod_1246(clk,rst,matrix_A[1246],matrix_B[46],mul_res1[1246]);
multi_7x28 multi_7x28_mod_1247(clk,rst,matrix_A[1247],matrix_B[47],mul_res1[1247]);
multi_7x28 multi_7x28_mod_1248(clk,rst,matrix_A[1248],matrix_B[48],mul_res1[1248]);
multi_7x28 multi_7x28_mod_1249(clk,rst,matrix_A[1249],matrix_B[49],mul_res1[1249]);
multi_7x28 multi_7x28_mod_1250(clk,rst,matrix_A[1250],matrix_B[50],mul_res1[1250]);
multi_7x28 multi_7x28_mod_1251(clk,rst,matrix_A[1251],matrix_B[51],mul_res1[1251]);
multi_7x28 multi_7x28_mod_1252(clk,rst,matrix_A[1252],matrix_B[52],mul_res1[1252]);
multi_7x28 multi_7x28_mod_1253(clk,rst,matrix_A[1253],matrix_B[53],mul_res1[1253]);
multi_7x28 multi_7x28_mod_1254(clk,rst,matrix_A[1254],matrix_B[54],mul_res1[1254]);
multi_7x28 multi_7x28_mod_1255(clk,rst,matrix_A[1255],matrix_B[55],mul_res1[1255]);
multi_7x28 multi_7x28_mod_1256(clk,rst,matrix_A[1256],matrix_B[56],mul_res1[1256]);
multi_7x28 multi_7x28_mod_1257(clk,rst,matrix_A[1257],matrix_B[57],mul_res1[1257]);
multi_7x28 multi_7x28_mod_1258(clk,rst,matrix_A[1258],matrix_B[58],mul_res1[1258]);
multi_7x28 multi_7x28_mod_1259(clk,rst,matrix_A[1259],matrix_B[59],mul_res1[1259]);
multi_7x28 multi_7x28_mod_1260(clk,rst,matrix_A[1260],matrix_B[60],mul_res1[1260]);
multi_7x28 multi_7x28_mod_1261(clk,rst,matrix_A[1261],matrix_B[61],mul_res1[1261]);
multi_7x28 multi_7x28_mod_1262(clk,rst,matrix_A[1262],matrix_B[62],mul_res1[1262]);
multi_7x28 multi_7x28_mod_1263(clk,rst,matrix_A[1263],matrix_B[63],mul_res1[1263]);
multi_7x28 multi_7x28_mod_1264(clk,rst,matrix_A[1264],matrix_B[64],mul_res1[1264]);
multi_7x28 multi_7x28_mod_1265(clk,rst,matrix_A[1265],matrix_B[65],mul_res1[1265]);
multi_7x28 multi_7x28_mod_1266(clk,rst,matrix_A[1266],matrix_B[66],mul_res1[1266]);
multi_7x28 multi_7x28_mod_1267(clk,rst,matrix_A[1267],matrix_B[67],mul_res1[1267]);
multi_7x28 multi_7x28_mod_1268(clk,rst,matrix_A[1268],matrix_B[68],mul_res1[1268]);
multi_7x28 multi_7x28_mod_1269(clk,rst,matrix_A[1269],matrix_B[69],mul_res1[1269]);
multi_7x28 multi_7x28_mod_1270(clk,rst,matrix_A[1270],matrix_B[70],mul_res1[1270]);
multi_7x28 multi_7x28_mod_1271(clk,rst,matrix_A[1271],matrix_B[71],mul_res1[1271]);
multi_7x28 multi_7x28_mod_1272(clk,rst,matrix_A[1272],matrix_B[72],mul_res1[1272]);
multi_7x28 multi_7x28_mod_1273(clk,rst,matrix_A[1273],matrix_B[73],mul_res1[1273]);
multi_7x28 multi_7x28_mod_1274(clk,rst,matrix_A[1274],matrix_B[74],mul_res1[1274]);
multi_7x28 multi_7x28_mod_1275(clk,rst,matrix_A[1275],matrix_B[75],mul_res1[1275]);
multi_7x28 multi_7x28_mod_1276(clk,rst,matrix_A[1276],matrix_B[76],mul_res1[1276]);
multi_7x28 multi_7x28_mod_1277(clk,rst,matrix_A[1277],matrix_B[77],mul_res1[1277]);
multi_7x28 multi_7x28_mod_1278(clk,rst,matrix_A[1278],matrix_B[78],mul_res1[1278]);
multi_7x28 multi_7x28_mod_1279(clk,rst,matrix_A[1279],matrix_B[79],mul_res1[1279]);
multi_7x28 multi_7x28_mod_1280(clk,rst,matrix_A[1280],matrix_B[80],mul_res1[1280]);
multi_7x28 multi_7x28_mod_1281(clk,rst,matrix_A[1281],matrix_B[81],mul_res1[1281]);
multi_7x28 multi_7x28_mod_1282(clk,rst,matrix_A[1282],matrix_B[82],mul_res1[1282]);
multi_7x28 multi_7x28_mod_1283(clk,rst,matrix_A[1283],matrix_B[83],mul_res1[1283]);
multi_7x28 multi_7x28_mod_1284(clk,rst,matrix_A[1284],matrix_B[84],mul_res1[1284]);
multi_7x28 multi_7x28_mod_1285(clk,rst,matrix_A[1285],matrix_B[85],mul_res1[1285]);
multi_7x28 multi_7x28_mod_1286(clk,rst,matrix_A[1286],matrix_B[86],mul_res1[1286]);
multi_7x28 multi_7x28_mod_1287(clk,rst,matrix_A[1287],matrix_B[87],mul_res1[1287]);
multi_7x28 multi_7x28_mod_1288(clk,rst,matrix_A[1288],matrix_B[88],mul_res1[1288]);
multi_7x28 multi_7x28_mod_1289(clk,rst,matrix_A[1289],matrix_B[89],mul_res1[1289]);
multi_7x28 multi_7x28_mod_1290(clk,rst,matrix_A[1290],matrix_B[90],mul_res1[1290]);
multi_7x28 multi_7x28_mod_1291(clk,rst,matrix_A[1291],matrix_B[91],mul_res1[1291]);
multi_7x28 multi_7x28_mod_1292(clk,rst,matrix_A[1292],matrix_B[92],mul_res1[1292]);
multi_7x28 multi_7x28_mod_1293(clk,rst,matrix_A[1293],matrix_B[93],mul_res1[1293]);
multi_7x28 multi_7x28_mod_1294(clk,rst,matrix_A[1294],matrix_B[94],mul_res1[1294]);
multi_7x28 multi_7x28_mod_1295(clk,rst,matrix_A[1295],matrix_B[95],mul_res1[1295]);
multi_7x28 multi_7x28_mod_1296(clk,rst,matrix_A[1296],matrix_B[96],mul_res1[1296]);
multi_7x28 multi_7x28_mod_1297(clk,rst,matrix_A[1297],matrix_B[97],mul_res1[1297]);
multi_7x28 multi_7x28_mod_1298(clk,rst,matrix_A[1298],matrix_B[98],mul_res1[1298]);
multi_7x28 multi_7x28_mod_1299(clk,rst,matrix_A[1299],matrix_B[99],mul_res1[1299]);
multi_7x28 multi_7x28_mod_1300(clk,rst,matrix_A[1300],matrix_B[100],mul_res1[1300]);
multi_7x28 multi_7x28_mod_1301(clk,rst,matrix_A[1301],matrix_B[101],mul_res1[1301]);
multi_7x28 multi_7x28_mod_1302(clk,rst,matrix_A[1302],matrix_B[102],mul_res1[1302]);
multi_7x28 multi_7x28_mod_1303(clk,rst,matrix_A[1303],matrix_B[103],mul_res1[1303]);
multi_7x28 multi_7x28_mod_1304(clk,rst,matrix_A[1304],matrix_B[104],mul_res1[1304]);
multi_7x28 multi_7x28_mod_1305(clk,rst,matrix_A[1305],matrix_B[105],mul_res1[1305]);
multi_7x28 multi_7x28_mod_1306(clk,rst,matrix_A[1306],matrix_B[106],mul_res1[1306]);
multi_7x28 multi_7x28_mod_1307(clk,rst,matrix_A[1307],matrix_B[107],mul_res1[1307]);
multi_7x28 multi_7x28_mod_1308(clk,rst,matrix_A[1308],matrix_B[108],mul_res1[1308]);
multi_7x28 multi_7x28_mod_1309(clk,rst,matrix_A[1309],matrix_B[109],mul_res1[1309]);
multi_7x28 multi_7x28_mod_1310(clk,rst,matrix_A[1310],matrix_B[110],mul_res1[1310]);
multi_7x28 multi_7x28_mod_1311(clk,rst,matrix_A[1311],matrix_B[111],mul_res1[1311]);
multi_7x28 multi_7x28_mod_1312(clk,rst,matrix_A[1312],matrix_B[112],mul_res1[1312]);
multi_7x28 multi_7x28_mod_1313(clk,rst,matrix_A[1313],matrix_B[113],mul_res1[1313]);
multi_7x28 multi_7x28_mod_1314(clk,rst,matrix_A[1314],matrix_B[114],mul_res1[1314]);
multi_7x28 multi_7x28_mod_1315(clk,rst,matrix_A[1315],matrix_B[115],mul_res1[1315]);
multi_7x28 multi_7x28_mod_1316(clk,rst,matrix_A[1316],matrix_B[116],mul_res1[1316]);
multi_7x28 multi_7x28_mod_1317(clk,rst,matrix_A[1317],matrix_B[117],mul_res1[1317]);
multi_7x28 multi_7x28_mod_1318(clk,rst,matrix_A[1318],matrix_B[118],mul_res1[1318]);
multi_7x28 multi_7x28_mod_1319(clk,rst,matrix_A[1319],matrix_B[119],mul_res1[1319]);
multi_7x28 multi_7x28_mod_1320(clk,rst,matrix_A[1320],matrix_B[120],mul_res1[1320]);
multi_7x28 multi_7x28_mod_1321(clk,rst,matrix_A[1321],matrix_B[121],mul_res1[1321]);
multi_7x28 multi_7x28_mod_1322(clk,rst,matrix_A[1322],matrix_B[122],mul_res1[1322]);
multi_7x28 multi_7x28_mod_1323(clk,rst,matrix_A[1323],matrix_B[123],mul_res1[1323]);
multi_7x28 multi_7x28_mod_1324(clk,rst,matrix_A[1324],matrix_B[124],mul_res1[1324]);
multi_7x28 multi_7x28_mod_1325(clk,rst,matrix_A[1325],matrix_B[125],mul_res1[1325]);
multi_7x28 multi_7x28_mod_1326(clk,rst,matrix_A[1326],matrix_B[126],mul_res1[1326]);
multi_7x28 multi_7x28_mod_1327(clk,rst,matrix_A[1327],matrix_B[127],mul_res1[1327]);
multi_7x28 multi_7x28_mod_1328(clk,rst,matrix_A[1328],matrix_B[128],mul_res1[1328]);
multi_7x28 multi_7x28_mod_1329(clk,rst,matrix_A[1329],matrix_B[129],mul_res1[1329]);
multi_7x28 multi_7x28_mod_1330(clk,rst,matrix_A[1330],matrix_B[130],mul_res1[1330]);
multi_7x28 multi_7x28_mod_1331(clk,rst,matrix_A[1331],matrix_B[131],mul_res1[1331]);
multi_7x28 multi_7x28_mod_1332(clk,rst,matrix_A[1332],matrix_B[132],mul_res1[1332]);
multi_7x28 multi_7x28_mod_1333(clk,rst,matrix_A[1333],matrix_B[133],mul_res1[1333]);
multi_7x28 multi_7x28_mod_1334(clk,rst,matrix_A[1334],matrix_B[134],mul_res1[1334]);
multi_7x28 multi_7x28_mod_1335(clk,rst,matrix_A[1335],matrix_B[135],mul_res1[1335]);
multi_7x28 multi_7x28_mod_1336(clk,rst,matrix_A[1336],matrix_B[136],mul_res1[1336]);
multi_7x28 multi_7x28_mod_1337(clk,rst,matrix_A[1337],matrix_B[137],mul_res1[1337]);
multi_7x28 multi_7x28_mod_1338(clk,rst,matrix_A[1338],matrix_B[138],mul_res1[1338]);
multi_7x28 multi_7x28_mod_1339(clk,rst,matrix_A[1339],matrix_B[139],mul_res1[1339]);
multi_7x28 multi_7x28_mod_1340(clk,rst,matrix_A[1340],matrix_B[140],mul_res1[1340]);
multi_7x28 multi_7x28_mod_1341(clk,rst,matrix_A[1341],matrix_B[141],mul_res1[1341]);
multi_7x28 multi_7x28_mod_1342(clk,rst,matrix_A[1342],matrix_B[142],mul_res1[1342]);
multi_7x28 multi_7x28_mod_1343(clk,rst,matrix_A[1343],matrix_B[143],mul_res1[1343]);
multi_7x28 multi_7x28_mod_1344(clk,rst,matrix_A[1344],matrix_B[144],mul_res1[1344]);
multi_7x28 multi_7x28_mod_1345(clk,rst,matrix_A[1345],matrix_B[145],mul_res1[1345]);
multi_7x28 multi_7x28_mod_1346(clk,rst,matrix_A[1346],matrix_B[146],mul_res1[1346]);
multi_7x28 multi_7x28_mod_1347(clk,rst,matrix_A[1347],matrix_B[147],mul_res1[1347]);
multi_7x28 multi_7x28_mod_1348(clk,rst,matrix_A[1348],matrix_B[148],mul_res1[1348]);
multi_7x28 multi_7x28_mod_1349(clk,rst,matrix_A[1349],matrix_B[149],mul_res1[1349]);
multi_7x28 multi_7x28_mod_1350(clk,rst,matrix_A[1350],matrix_B[150],mul_res1[1350]);
multi_7x28 multi_7x28_mod_1351(clk,rst,matrix_A[1351],matrix_B[151],mul_res1[1351]);
multi_7x28 multi_7x28_mod_1352(clk,rst,matrix_A[1352],matrix_B[152],mul_res1[1352]);
multi_7x28 multi_7x28_mod_1353(clk,rst,matrix_A[1353],matrix_B[153],mul_res1[1353]);
multi_7x28 multi_7x28_mod_1354(clk,rst,matrix_A[1354],matrix_B[154],mul_res1[1354]);
multi_7x28 multi_7x28_mod_1355(clk,rst,matrix_A[1355],matrix_B[155],mul_res1[1355]);
multi_7x28 multi_7x28_mod_1356(clk,rst,matrix_A[1356],matrix_B[156],mul_res1[1356]);
multi_7x28 multi_7x28_mod_1357(clk,rst,matrix_A[1357],matrix_B[157],mul_res1[1357]);
multi_7x28 multi_7x28_mod_1358(clk,rst,matrix_A[1358],matrix_B[158],mul_res1[1358]);
multi_7x28 multi_7x28_mod_1359(clk,rst,matrix_A[1359],matrix_B[159],mul_res1[1359]);
multi_7x28 multi_7x28_mod_1360(clk,rst,matrix_A[1360],matrix_B[160],mul_res1[1360]);
multi_7x28 multi_7x28_mod_1361(clk,rst,matrix_A[1361],matrix_B[161],mul_res1[1361]);
multi_7x28 multi_7x28_mod_1362(clk,rst,matrix_A[1362],matrix_B[162],mul_res1[1362]);
multi_7x28 multi_7x28_mod_1363(clk,rst,matrix_A[1363],matrix_B[163],mul_res1[1363]);
multi_7x28 multi_7x28_mod_1364(clk,rst,matrix_A[1364],matrix_B[164],mul_res1[1364]);
multi_7x28 multi_7x28_mod_1365(clk,rst,matrix_A[1365],matrix_B[165],mul_res1[1365]);
multi_7x28 multi_7x28_mod_1366(clk,rst,matrix_A[1366],matrix_B[166],mul_res1[1366]);
multi_7x28 multi_7x28_mod_1367(clk,rst,matrix_A[1367],matrix_B[167],mul_res1[1367]);
multi_7x28 multi_7x28_mod_1368(clk,rst,matrix_A[1368],matrix_B[168],mul_res1[1368]);
multi_7x28 multi_7x28_mod_1369(clk,rst,matrix_A[1369],matrix_B[169],mul_res1[1369]);
multi_7x28 multi_7x28_mod_1370(clk,rst,matrix_A[1370],matrix_B[170],mul_res1[1370]);
multi_7x28 multi_7x28_mod_1371(clk,rst,matrix_A[1371],matrix_B[171],mul_res1[1371]);
multi_7x28 multi_7x28_mod_1372(clk,rst,matrix_A[1372],matrix_B[172],mul_res1[1372]);
multi_7x28 multi_7x28_mod_1373(clk,rst,matrix_A[1373],matrix_B[173],mul_res1[1373]);
multi_7x28 multi_7x28_mod_1374(clk,rst,matrix_A[1374],matrix_B[174],mul_res1[1374]);
multi_7x28 multi_7x28_mod_1375(clk,rst,matrix_A[1375],matrix_B[175],mul_res1[1375]);
multi_7x28 multi_7x28_mod_1376(clk,rst,matrix_A[1376],matrix_B[176],mul_res1[1376]);
multi_7x28 multi_7x28_mod_1377(clk,rst,matrix_A[1377],matrix_B[177],mul_res1[1377]);
multi_7x28 multi_7x28_mod_1378(clk,rst,matrix_A[1378],matrix_B[178],mul_res1[1378]);
multi_7x28 multi_7x28_mod_1379(clk,rst,matrix_A[1379],matrix_B[179],mul_res1[1379]);
multi_7x28 multi_7x28_mod_1380(clk,rst,matrix_A[1380],matrix_B[180],mul_res1[1380]);
multi_7x28 multi_7x28_mod_1381(clk,rst,matrix_A[1381],matrix_B[181],mul_res1[1381]);
multi_7x28 multi_7x28_mod_1382(clk,rst,matrix_A[1382],matrix_B[182],mul_res1[1382]);
multi_7x28 multi_7x28_mod_1383(clk,rst,matrix_A[1383],matrix_B[183],mul_res1[1383]);
multi_7x28 multi_7x28_mod_1384(clk,rst,matrix_A[1384],matrix_B[184],mul_res1[1384]);
multi_7x28 multi_7x28_mod_1385(clk,rst,matrix_A[1385],matrix_B[185],mul_res1[1385]);
multi_7x28 multi_7x28_mod_1386(clk,rst,matrix_A[1386],matrix_B[186],mul_res1[1386]);
multi_7x28 multi_7x28_mod_1387(clk,rst,matrix_A[1387],matrix_B[187],mul_res1[1387]);
multi_7x28 multi_7x28_mod_1388(clk,rst,matrix_A[1388],matrix_B[188],mul_res1[1388]);
multi_7x28 multi_7x28_mod_1389(clk,rst,matrix_A[1389],matrix_B[189],mul_res1[1389]);
multi_7x28 multi_7x28_mod_1390(clk,rst,matrix_A[1390],matrix_B[190],mul_res1[1390]);
multi_7x28 multi_7x28_mod_1391(clk,rst,matrix_A[1391],matrix_B[191],mul_res1[1391]);
multi_7x28 multi_7x28_mod_1392(clk,rst,matrix_A[1392],matrix_B[192],mul_res1[1392]);
multi_7x28 multi_7x28_mod_1393(clk,rst,matrix_A[1393],matrix_B[193],mul_res1[1393]);
multi_7x28 multi_7x28_mod_1394(clk,rst,matrix_A[1394],matrix_B[194],mul_res1[1394]);
multi_7x28 multi_7x28_mod_1395(clk,rst,matrix_A[1395],matrix_B[195],mul_res1[1395]);
multi_7x28 multi_7x28_mod_1396(clk,rst,matrix_A[1396],matrix_B[196],mul_res1[1396]);
multi_7x28 multi_7x28_mod_1397(clk,rst,matrix_A[1397],matrix_B[197],mul_res1[1397]);
multi_7x28 multi_7x28_mod_1398(clk,rst,matrix_A[1398],matrix_B[198],mul_res1[1398]);
multi_7x28 multi_7x28_mod_1399(clk,rst,matrix_A[1399],matrix_B[199],mul_res1[1399]);
multi_7x28 multi_7x28_mod_1400(clk,rst,matrix_A[1400],matrix_B[0],mul_res1[1400]);
multi_7x28 multi_7x28_mod_1401(clk,rst,matrix_A[1401],matrix_B[1],mul_res1[1401]);
multi_7x28 multi_7x28_mod_1402(clk,rst,matrix_A[1402],matrix_B[2],mul_res1[1402]);
multi_7x28 multi_7x28_mod_1403(clk,rst,matrix_A[1403],matrix_B[3],mul_res1[1403]);
multi_7x28 multi_7x28_mod_1404(clk,rst,matrix_A[1404],matrix_B[4],mul_res1[1404]);
multi_7x28 multi_7x28_mod_1405(clk,rst,matrix_A[1405],matrix_B[5],mul_res1[1405]);
multi_7x28 multi_7x28_mod_1406(clk,rst,matrix_A[1406],matrix_B[6],mul_res1[1406]);
multi_7x28 multi_7x28_mod_1407(clk,rst,matrix_A[1407],matrix_B[7],mul_res1[1407]);
multi_7x28 multi_7x28_mod_1408(clk,rst,matrix_A[1408],matrix_B[8],mul_res1[1408]);
multi_7x28 multi_7x28_mod_1409(clk,rst,matrix_A[1409],matrix_B[9],mul_res1[1409]);
multi_7x28 multi_7x28_mod_1410(clk,rst,matrix_A[1410],matrix_B[10],mul_res1[1410]);
multi_7x28 multi_7x28_mod_1411(clk,rst,matrix_A[1411],matrix_B[11],mul_res1[1411]);
multi_7x28 multi_7x28_mod_1412(clk,rst,matrix_A[1412],matrix_B[12],mul_res1[1412]);
multi_7x28 multi_7x28_mod_1413(clk,rst,matrix_A[1413],matrix_B[13],mul_res1[1413]);
multi_7x28 multi_7x28_mod_1414(clk,rst,matrix_A[1414],matrix_B[14],mul_res1[1414]);
multi_7x28 multi_7x28_mod_1415(clk,rst,matrix_A[1415],matrix_B[15],mul_res1[1415]);
multi_7x28 multi_7x28_mod_1416(clk,rst,matrix_A[1416],matrix_B[16],mul_res1[1416]);
multi_7x28 multi_7x28_mod_1417(clk,rst,matrix_A[1417],matrix_B[17],mul_res1[1417]);
multi_7x28 multi_7x28_mod_1418(clk,rst,matrix_A[1418],matrix_B[18],mul_res1[1418]);
multi_7x28 multi_7x28_mod_1419(clk,rst,matrix_A[1419],matrix_B[19],mul_res1[1419]);
multi_7x28 multi_7x28_mod_1420(clk,rst,matrix_A[1420],matrix_B[20],mul_res1[1420]);
multi_7x28 multi_7x28_mod_1421(clk,rst,matrix_A[1421],matrix_B[21],mul_res1[1421]);
multi_7x28 multi_7x28_mod_1422(clk,rst,matrix_A[1422],matrix_B[22],mul_res1[1422]);
multi_7x28 multi_7x28_mod_1423(clk,rst,matrix_A[1423],matrix_B[23],mul_res1[1423]);
multi_7x28 multi_7x28_mod_1424(clk,rst,matrix_A[1424],matrix_B[24],mul_res1[1424]);
multi_7x28 multi_7x28_mod_1425(clk,rst,matrix_A[1425],matrix_B[25],mul_res1[1425]);
multi_7x28 multi_7x28_mod_1426(clk,rst,matrix_A[1426],matrix_B[26],mul_res1[1426]);
multi_7x28 multi_7x28_mod_1427(clk,rst,matrix_A[1427],matrix_B[27],mul_res1[1427]);
multi_7x28 multi_7x28_mod_1428(clk,rst,matrix_A[1428],matrix_B[28],mul_res1[1428]);
multi_7x28 multi_7x28_mod_1429(clk,rst,matrix_A[1429],matrix_B[29],mul_res1[1429]);
multi_7x28 multi_7x28_mod_1430(clk,rst,matrix_A[1430],matrix_B[30],mul_res1[1430]);
multi_7x28 multi_7x28_mod_1431(clk,rst,matrix_A[1431],matrix_B[31],mul_res1[1431]);
multi_7x28 multi_7x28_mod_1432(clk,rst,matrix_A[1432],matrix_B[32],mul_res1[1432]);
multi_7x28 multi_7x28_mod_1433(clk,rst,matrix_A[1433],matrix_B[33],mul_res1[1433]);
multi_7x28 multi_7x28_mod_1434(clk,rst,matrix_A[1434],matrix_B[34],mul_res1[1434]);
multi_7x28 multi_7x28_mod_1435(clk,rst,matrix_A[1435],matrix_B[35],mul_res1[1435]);
multi_7x28 multi_7x28_mod_1436(clk,rst,matrix_A[1436],matrix_B[36],mul_res1[1436]);
multi_7x28 multi_7x28_mod_1437(clk,rst,matrix_A[1437],matrix_B[37],mul_res1[1437]);
multi_7x28 multi_7x28_mod_1438(clk,rst,matrix_A[1438],matrix_B[38],mul_res1[1438]);
multi_7x28 multi_7x28_mod_1439(clk,rst,matrix_A[1439],matrix_B[39],mul_res1[1439]);
multi_7x28 multi_7x28_mod_1440(clk,rst,matrix_A[1440],matrix_B[40],mul_res1[1440]);
multi_7x28 multi_7x28_mod_1441(clk,rst,matrix_A[1441],matrix_B[41],mul_res1[1441]);
multi_7x28 multi_7x28_mod_1442(clk,rst,matrix_A[1442],matrix_B[42],mul_res1[1442]);
multi_7x28 multi_7x28_mod_1443(clk,rst,matrix_A[1443],matrix_B[43],mul_res1[1443]);
multi_7x28 multi_7x28_mod_1444(clk,rst,matrix_A[1444],matrix_B[44],mul_res1[1444]);
multi_7x28 multi_7x28_mod_1445(clk,rst,matrix_A[1445],matrix_B[45],mul_res1[1445]);
multi_7x28 multi_7x28_mod_1446(clk,rst,matrix_A[1446],matrix_B[46],mul_res1[1446]);
multi_7x28 multi_7x28_mod_1447(clk,rst,matrix_A[1447],matrix_B[47],mul_res1[1447]);
multi_7x28 multi_7x28_mod_1448(clk,rst,matrix_A[1448],matrix_B[48],mul_res1[1448]);
multi_7x28 multi_7x28_mod_1449(clk,rst,matrix_A[1449],matrix_B[49],mul_res1[1449]);
multi_7x28 multi_7x28_mod_1450(clk,rst,matrix_A[1450],matrix_B[50],mul_res1[1450]);
multi_7x28 multi_7x28_mod_1451(clk,rst,matrix_A[1451],matrix_B[51],mul_res1[1451]);
multi_7x28 multi_7x28_mod_1452(clk,rst,matrix_A[1452],matrix_B[52],mul_res1[1452]);
multi_7x28 multi_7x28_mod_1453(clk,rst,matrix_A[1453],matrix_B[53],mul_res1[1453]);
multi_7x28 multi_7x28_mod_1454(clk,rst,matrix_A[1454],matrix_B[54],mul_res1[1454]);
multi_7x28 multi_7x28_mod_1455(clk,rst,matrix_A[1455],matrix_B[55],mul_res1[1455]);
multi_7x28 multi_7x28_mod_1456(clk,rst,matrix_A[1456],matrix_B[56],mul_res1[1456]);
multi_7x28 multi_7x28_mod_1457(clk,rst,matrix_A[1457],matrix_B[57],mul_res1[1457]);
multi_7x28 multi_7x28_mod_1458(clk,rst,matrix_A[1458],matrix_B[58],mul_res1[1458]);
multi_7x28 multi_7x28_mod_1459(clk,rst,matrix_A[1459],matrix_B[59],mul_res1[1459]);
multi_7x28 multi_7x28_mod_1460(clk,rst,matrix_A[1460],matrix_B[60],mul_res1[1460]);
multi_7x28 multi_7x28_mod_1461(clk,rst,matrix_A[1461],matrix_B[61],mul_res1[1461]);
multi_7x28 multi_7x28_mod_1462(clk,rst,matrix_A[1462],matrix_B[62],mul_res1[1462]);
multi_7x28 multi_7x28_mod_1463(clk,rst,matrix_A[1463],matrix_B[63],mul_res1[1463]);
multi_7x28 multi_7x28_mod_1464(clk,rst,matrix_A[1464],matrix_B[64],mul_res1[1464]);
multi_7x28 multi_7x28_mod_1465(clk,rst,matrix_A[1465],matrix_B[65],mul_res1[1465]);
multi_7x28 multi_7x28_mod_1466(clk,rst,matrix_A[1466],matrix_B[66],mul_res1[1466]);
multi_7x28 multi_7x28_mod_1467(clk,rst,matrix_A[1467],matrix_B[67],mul_res1[1467]);
multi_7x28 multi_7x28_mod_1468(clk,rst,matrix_A[1468],matrix_B[68],mul_res1[1468]);
multi_7x28 multi_7x28_mod_1469(clk,rst,matrix_A[1469],matrix_B[69],mul_res1[1469]);
multi_7x28 multi_7x28_mod_1470(clk,rst,matrix_A[1470],matrix_B[70],mul_res1[1470]);
multi_7x28 multi_7x28_mod_1471(clk,rst,matrix_A[1471],matrix_B[71],mul_res1[1471]);
multi_7x28 multi_7x28_mod_1472(clk,rst,matrix_A[1472],matrix_B[72],mul_res1[1472]);
multi_7x28 multi_7x28_mod_1473(clk,rst,matrix_A[1473],matrix_B[73],mul_res1[1473]);
multi_7x28 multi_7x28_mod_1474(clk,rst,matrix_A[1474],matrix_B[74],mul_res1[1474]);
multi_7x28 multi_7x28_mod_1475(clk,rst,matrix_A[1475],matrix_B[75],mul_res1[1475]);
multi_7x28 multi_7x28_mod_1476(clk,rst,matrix_A[1476],matrix_B[76],mul_res1[1476]);
multi_7x28 multi_7x28_mod_1477(clk,rst,matrix_A[1477],matrix_B[77],mul_res1[1477]);
multi_7x28 multi_7x28_mod_1478(clk,rst,matrix_A[1478],matrix_B[78],mul_res1[1478]);
multi_7x28 multi_7x28_mod_1479(clk,rst,matrix_A[1479],matrix_B[79],mul_res1[1479]);
multi_7x28 multi_7x28_mod_1480(clk,rst,matrix_A[1480],matrix_B[80],mul_res1[1480]);
multi_7x28 multi_7x28_mod_1481(clk,rst,matrix_A[1481],matrix_B[81],mul_res1[1481]);
multi_7x28 multi_7x28_mod_1482(clk,rst,matrix_A[1482],matrix_B[82],mul_res1[1482]);
multi_7x28 multi_7x28_mod_1483(clk,rst,matrix_A[1483],matrix_B[83],mul_res1[1483]);
multi_7x28 multi_7x28_mod_1484(clk,rst,matrix_A[1484],matrix_B[84],mul_res1[1484]);
multi_7x28 multi_7x28_mod_1485(clk,rst,matrix_A[1485],matrix_B[85],mul_res1[1485]);
multi_7x28 multi_7x28_mod_1486(clk,rst,matrix_A[1486],matrix_B[86],mul_res1[1486]);
multi_7x28 multi_7x28_mod_1487(clk,rst,matrix_A[1487],matrix_B[87],mul_res1[1487]);
multi_7x28 multi_7x28_mod_1488(clk,rst,matrix_A[1488],matrix_B[88],mul_res1[1488]);
multi_7x28 multi_7x28_mod_1489(clk,rst,matrix_A[1489],matrix_B[89],mul_res1[1489]);
multi_7x28 multi_7x28_mod_1490(clk,rst,matrix_A[1490],matrix_B[90],mul_res1[1490]);
multi_7x28 multi_7x28_mod_1491(clk,rst,matrix_A[1491],matrix_B[91],mul_res1[1491]);
multi_7x28 multi_7x28_mod_1492(clk,rst,matrix_A[1492],matrix_B[92],mul_res1[1492]);
multi_7x28 multi_7x28_mod_1493(clk,rst,matrix_A[1493],matrix_B[93],mul_res1[1493]);
multi_7x28 multi_7x28_mod_1494(clk,rst,matrix_A[1494],matrix_B[94],mul_res1[1494]);
multi_7x28 multi_7x28_mod_1495(clk,rst,matrix_A[1495],matrix_B[95],mul_res1[1495]);
multi_7x28 multi_7x28_mod_1496(clk,rst,matrix_A[1496],matrix_B[96],mul_res1[1496]);
multi_7x28 multi_7x28_mod_1497(clk,rst,matrix_A[1497],matrix_B[97],mul_res1[1497]);
multi_7x28 multi_7x28_mod_1498(clk,rst,matrix_A[1498],matrix_B[98],mul_res1[1498]);
multi_7x28 multi_7x28_mod_1499(clk,rst,matrix_A[1499],matrix_B[99],mul_res1[1499]);
multi_7x28 multi_7x28_mod_1500(clk,rst,matrix_A[1500],matrix_B[100],mul_res1[1500]);
multi_7x28 multi_7x28_mod_1501(clk,rst,matrix_A[1501],matrix_B[101],mul_res1[1501]);
multi_7x28 multi_7x28_mod_1502(clk,rst,matrix_A[1502],matrix_B[102],mul_res1[1502]);
multi_7x28 multi_7x28_mod_1503(clk,rst,matrix_A[1503],matrix_B[103],mul_res1[1503]);
multi_7x28 multi_7x28_mod_1504(clk,rst,matrix_A[1504],matrix_B[104],mul_res1[1504]);
multi_7x28 multi_7x28_mod_1505(clk,rst,matrix_A[1505],matrix_B[105],mul_res1[1505]);
multi_7x28 multi_7x28_mod_1506(clk,rst,matrix_A[1506],matrix_B[106],mul_res1[1506]);
multi_7x28 multi_7x28_mod_1507(clk,rst,matrix_A[1507],matrix_B[107],mul_res1[1507]);
multi_7x28 multi_7x28_mod_1508(clk,rst,matrix_A[1508],matrix_B[108],mul_res1[1508]);
multi_7x28 multi_7x28_mod_1509(clk,rst,matrix_A[1509],matrix_B[109],mul_res1[1509]);
multi_7x28 multi_7x28_mod_1510(clk,rst,matrix_A[1510],matrix_B[110],mul_res1[1510]);
multi_7x28 multi_7x28_mod_1511(clk,rst,matrix_A[1511],matrix_B[111],mul_res1[1511]);
multi_7x28 multi_7x28_mod_1512(clk,rst,matrix_A[1512],matrix_B[112],mul_res1[1512]);
multi_7x28 multi_7x28_mod_1513(clk,rst,matrix_A[1513],matrix_B[113],mul_res1[1513]);
multi_7x28 multi_7x28_mod_1514(clk,rst,matrix_A[1514],matrix_B[114],mul_res1[1514]);
multi_7x28 multi_7x28_mod_1515(clk,rst,matrix_A[1515],matrix_B[115],mul_res1[1515]);
multi_7x28 multi_7x28_mod_1516(clk,rst,matrix_A[1516],matrix_B[116],mul_res1[1516]);
multi_7x28 multi_7x28_mod_1517(clk,rst,matrix_A[1517],matrix_B[117],mul_res1[1517]);
multi_7x28 multi_7x28_mod_1518(clk,rst,matrix_A[1518],matrix_B[118],mul_res1[1518]);
multi_7x28 multi_7x28_mod_1519(clk,rst,matrix_A[1519],matrix_B[119],mul_res1[1519]);
multi_7x28 multi_7x28_mod_1520(clk,rst,matrix_A[1520],matrix_B[120],mul_res1[1520]);
multi_7x28 multi_7x28_mod_1521(clk,rst,matrix_A[1521],matrix_B[121],mul_res1[1521]);
multi_7x28 multi_7x28_mod_1522(clk,rst,matrix_A[1522],matrix_B[122],mul_res1[1522]);
multi_7x28 multi_7x28_mod_1523(clk,rst,matrix_A[1523],matrix_B[123],mul_res1[1523]);
multi_7x28 multi_7x28_mod_1524(clk,rst,matrix_A[1524],matrix_B[124],mul_res1[1524]);
multi_7x28 multi_7x28_mod_1525(clk,rst,matrix_A[1525],matrix_B[125],mul_res1[1525]);
multi_7x28 multi_7x28_mod_1526(clk,rst,matrix_A[1526],matrix_B[126],mul_res1[1526]);
multi_7x28 multi_7x28_mod_1527(clk,rst,matrix_A[1527],matrix_B[127],mul_res1[1527]);
multi_7x28 multi_7x28_mod_1528(clk,rst,matrix_A[1528],matrix_B[128],mul_res1[1528]);
multi_7x28 multi_7x28_mod_1529(clk,rst,matrix_A[1529],matrix_B[129],mul_res1[1529]);
multi_7x28 multi_7x28_mod_1530(clk,rst,matrix_A[1530],matrix_B[130],mul_res1[1530]);
multi_7x28 multi_7x28_mod_1531(clk,rst,matrix_A[1531],matrix_B[131],mul_res1[1531]);
multi_7x28 multi_7x28_mod_1532(clk,rst,matrix_A[1532],matrix_B[132],mul_res1[1532]);
multi_7x28 multi_7x28_mod_1533(clk,rst,matrix_A[1533],matrix_B[133],mul_res1[1533]);
multi_7x28 multi_7x28_mod_1534(clk,rst,matrix_A[1534],matrix_B[134],mul_res1[1534]);
multi_7x28 multi_7x28_mod_1535(clk,rst,matrix_A[1535],matrix_B[135],mul_res1[1535]);
multi_7x28 multi_7x28_mod_1536(clk,rst,matrix_A[1536],matrix_B[136],mul_res1[1536]);
multi_7x28 multi_7x28_mod_1537(clk,rst,matrix_A[1537],matrix_B[137],mul_res1[1537]);
multi_7x28 multi_7x28_mod_1538(clk,rst,matrix_A[1538],matrix_B[138],mul_res1[1538]);
multi_7x28 multi_7x28_mod_1539(clk,rst,matrix_A[1539],matrix_B[139],mul_res1[1539]);
multi_7x28 multi_7x28_mod_1540(clk,rst,matrix_A[1540],matrix_B[140],mul_res1[1540]);
multi_7x28 multi_7x28_mod_1541(clk,rst,matrix_A[1541],matrix_B[141],mul_res1[1541]);
multi_7x28 multi_7x28_mod_1542(clk,rst,matrix_A[1542],matrix_B[142],mul_res1[1542]);
multi_7x28 multi_7x28_mod_1543(clk,rst,matrix_A[1543],matrix_B[143],mul_res1[1543]);
multi_7x28 multi_7x28_mod_1544(clk,rst,matrix_A[1544],matrix_B[144],mul_res1[1544]);
multi_7x28 multi_7x28_mod_1545(clk,rst,matrix_A[1545],matrix_B[145],mul_res1[1545]);
multi_7x28 multi_7x28_mod_1546(clk,rst,matrix_A[1546],matrix_B[146],mul_res1[1546]);
multi_7x28 multi_7x28_mod_1547(clk,rst,matrix_A[1547],matrix_B[147],mul_res1[1547]);
multi_7x28 multi_7x28_mod_1548(clk,rst,matrix_A[1548],matrix_B[148],mul_res1[1548]);
multi_7x28 multi_7x28_mod_1549(clk,rst,matrix_A[1549],matrix_B[149],mul_res1[1549]);
multi_7x28 multi_7x28_mod_1550(clk,rst,matrix_A[1550],matrix_B[150],mul_res1[1550]);
multi_7x28 multi_7x28_mod_1551(clk,rst,matrix_A[1551],matrix_B[151],mul_res1[1551]);
multi_7x28 multi_7x28_mod_1552(clk,rst,matrix_A[1552],matrix_B[152],mul_res1[1552]);
multi_7x28 multi_7x28_mod_1553(clk,rst,matrix_A[1553],matrix_B[153],mul_res1[1553]);
multi_7x28 multi_7x28_mod_1554(clk,rst,matrix_A[1554],matrix_B[154],mul_res1[1554]);
multi_7x28 multi_7x28_mod_1555(clk,rst,matrix_A[1555],matrix_B[155],mul_res1[1555]);
multi_7x28 multi_7x28_mod_1556(clk,rst,matrix_A[1556],matrix_B[156],mul_res1[1556]);
multi_7x28 multi_7x28_mod_1557(clk,rst,matrix_A[1557],matrix_B[157],mul_res1[1557]);
multi_7x28 multi_7x28_mod_1558(clk,rst,matrix_A[1558],matrix_B[158],mul_res1[1558]);
multi_7x28 multi_7x28_mod_1559(clk,rst,matrix_A[1559],matrix_B[159],mul_res1[1559]);
multi_7x28 multi_7x28_mod_1560(clk,rst,matrix_A[1560],matrix_B[160],mul_res1[1560]);
multi_7x28 multi_7x28_mod_1561(clk,rst,matrix_A[1561],matrix_B[161],mul_res1[1561]);
multi_7x28 multi_7x28_mod_1562(clk,rst,matrix_A[1562],matrix_B[162],mul_res1[1562]);
multi_7x28 multi_7x28_mod_1563(clk,rst,matrix_A[1563],matrix_B[163],mul_res1[1563]);
multi_7x28 multi_7x28_mod_1564(clk,rst,matrix_A[1564],matrix_B[164],mul_res1[1564]);
multi_7x28 multi_7x28_mod_1565(clk,rst,matrix_A[1565],matrix_B[165],mul_res1[1565]);
multi_7x28 multi_7x28_mod_1566(clk,rst,matrix_A[1566],matrix_B[166],mul_res1[1566]);
multi_7x28 multi_7x28_mod_1567(clk,rst,matrix_A[1567],matrix_B[167],mul_res1[1567]);
multi_7x28 multi_7x28_mod_1568(clk,rst,matrix_A[1568],matrix_B[168],mul_res1[1568]);
multi_7x28 multi_7x28_mod_1569(clk,rst,matrix_A[1569],matrix_B[169],mul_res1[1569]);
multi_7x28 multi_7x28_mod_1570(clk,rst,matrix_A[1570],matrix_B[170],mul_res1[1570]);
multi_7x28 multi_7x28_mod_1571(clk,rst,matrix_A[1571],matrix_B[171],mul_res1[1571]);
multi_7x28 multi_7x28_mod_1572(clk,rst,matrix_A[1572],matrix_B[172],mul_res1[1572]);
multi_7x28 multi_7x28_mod_1573(clk,rst,matrix_A[1573],matrix_B[173],mul_res1[1573]);
multi_7x28 multi_7x28_mod_1574(clk,rst,matrix_A[1574],matrix_B[174],mul_res1[1574]);
multi_7x28 multi_7x28_mod_1575(clk,rst,matrix_A[1575],matrix_B[175],mul_res1[1575]);
multi_7x28 multi_7x28_mod_1576(clk,rst,matrix_A[1576],matrix_B[176],mul_res1[1576]);
multi_7x28 multi_7x28_mod_1577(clk,rst,matrix_A[1577],matrix_B[177],mul_res1[1577]);
multi_7x28 multi_7x28_mod_1578(clk,rst,matrix_A[1578],matrix_B[178],mul_res1[1578]);
multi_7x28 multi_7x28_mod_1579(clk,rst,matrix_A[1579],matrix_B[179],mul_res1[1579]);
multi_7x28 multi_7x28_mod_1580(clk,rst,matrix_A[1580],matrix_B[180],mul_res1[1580]);
multi_7x28 multi_7x28_mod_1581(clk,rst,matrix_A[1581],matrix_B[181],mul_res1[1581]);
multi_7x28 multi_7x28_mod_1582(clk,rst,matrix_A[1582],matrix_B[182],mul_res1[1582]);
multi_7x28 multi_7x28_mod_1583(clk,rst,matrix_A[1583],matrix_B[183],mul_res1[1583]);
multi_7x28 multi_7x28_mod_1584(clk,rst,matrix_A[1584],matrix_B[184],mul_res1[1584]);
multi_7x28 multi_7x28_mod_1585(clk,rst,matrix_A[1585],matrix_B[185],mul_res1[1585]);
multi_7x28 multi_7x28_mod_1586(clk,rst,matrix_A[1586],matrix_B[186],mul_res1[1586]);
multi_7x28 multi_7x28_mod_1587(clk,rst,matrix_A[1587],matrix_B[187],mul_res1[1587]);
multi_7x28 multi_7x28_mod_1588(clk,rst,matrix_A[1588],matrix_B[188],mul_res1[1588]);
multi_7x28 multi_7x28_mod_1589(clk,rst,matrix_A[1589],matrix_B[189],mul_res1[1589]);
multi_7x28 multi_7x28_mod_1590(clk,rst,matrix_A[1590],matrix_B[190],mul_res1[1590]);
multi_7x28 multi_7x28_mod_1591(clk,rst,matrix_A[1591],matrix_B[191],mul_res1[1591]);
multi_7x28 multi_7x28_mod_1592(clk,rst,matrix_A[1592],matrix_B[192],mul_res1[1592]);
multi_7x28 multi_7x28_mod_1593(clk,rst,matrix_A[1593],matrix_B[193],mul_res1[1593]);
multi_7x28 multi_7x28_mod_1594(clk,rst,matrix_A[1594],matrix_B[194],mul_res1[1594]);
multi_7x28 multi_7x28_mod_1595(clk,rst,matrix_A[1595],matrix_B[195],mul_res1[1595]);
multi_7x28 multi_7x28_mod_1596(clk,rst,matrix_A[1596],matrix_B[196],mul_res1[1596]);
multi_7x28 multi_7x28_mod_1597(clk,rst,matrix_A[1597],matrix_B[197],mul_res1[1597]);
multi_7x28 multi_7x28_mod_1598(clk,rst,matrix_A[1598],matrix_B[198],mul_res1[1598]);
multi_7x28 multi_7x28_mod_1599(clk,rst,matrix_A[1599],matrix_B[199],mul_res1[1599]);
multi_7x28 multi_7x28_mod_1600(clk,rst,matrix_A[1600],matrix_B[0],mul_res1[1600]);
multi_7x28 multi_7x28_mod_1601(clk,rst,matrix_A[1601],matrix_B[1],mul_res1[1601]);
multi_7x28 multi_7x28_mod_1602(clk,rst,matrix_A[1602],matrix_B[2],mul_res1[1602]);
multi_7x28 multi_7x28_mod_1603(clk,rst,matrix_A[1603],matrix_B[3],mul_res1[1603]);
multi_7x28 multi_7x28_mod_1604(clk,rst,matrix_A[1604],matrix_B[4],mul_res1[1604]);
multi_7x28 multi_7x28_mod_1605(clk,rst,matrix_A[1605],matrix_B[5],mul_res1[1605]);
multi_7x28 multi_7x28_mod_1606(clk,rst,matrix_A[1606],matrix_B[6],mul_res1[1606]);
multi_7x28 multi_7x28_mod_1607(clk,rst,matrix_A[1607],matrix_B[7],mul_res1[1607]);
multi_7x28 multi_7x28_mod_1608(clk,rst,matrix_A[1608],matrix_B[8],mul_res1[1608]);
multi_7x28 multi_7x28_mod_1609(clk,rst,matrix_A[1609],matrix_B[9],mul_res1[1609]);
multi_7x28 multi_7x28_mod_1610(clk,rst,matrix_A[1610],matrix_B[10],mul_res1[1610]);
multi_7x28 multi_7x28_mod_1611(clk,rst,matrix_A[1611],matrix_B[11],mul_res1[1611]);
multi_7x28 multi_7x28_mod_1612(clk,rst,matrix_A[1612],matrix_B[12],mul_res1[1612]);
multi_7x28 multi_7x28_mod_1613(clk,rst,matrix_A[1613],matrix_B[13],mul_res1[1613]);
multi_7x28 multi_7x28_mod_1614(clk,rst,matrix_A[1614],matrix_B[14],mul_res1[1614]);
multi_7x28 multi_7x28_mod_1615(clk,rst,matrix_A[1615],matrix_B[15],mul_res1[1615]);
multi_7x28 multi_7x28_mod_1616(clk,rst,matrix_A[1616],matrix_B[16],mul_res1[1616]);
multi_7x28 multi_7x28_mod_1617(clk,rst,matrix_A[1617],matrix_B[17],mul_res1[1617]);
multi_7x28 multi_7x28_mod_1618(clk,rst,matrix_A[1618],matrix_B[18],mul_res1[1618]);
multi_7x28 multi_7x28_mod_1619(clk,rst,matrix_A[1619],matrix_B[19],mul_res1[1619]);
multi_7x28 multi_7x28_mod_1620(clk,rst,matrix_A[1620],matrix_B[20],mul_res1[1620]);
multi_7x28 multi_7x28_mod_1621(clk,rst,matrix_A[1621],matrix_B[21],mul_res1[1621]);
multi_7x28 multi_7x28_mod_1622(clk,rst,matrix_A[1622],matrix_B[22],mul_res1[1622]);
multi_7x28 multi_7x28_mod_1623(clk,rst,matrix_A[1623],matrix_B[23],mul_res1[1623]);
multi_7x28 multi_7x28_mod_1624(clk,rst,matrix_A[1624],matrix_B[24],mul_res1[1624]);
multi_7x28 multi_7x28_mod_1625(clk,rst,matrix_A[1625],matrix_B[25],mul_res1[1625]);
multi_7x28 multi_7x28_mod_1626(clk,rst,matrix_A[1626],matrix_B[26],mul_res1[1626]);
multi_7x28 multi_7x28_mod_1627(clk,rst,matrix_A[1627],matrix_B[27],mul_res1[1627]);
multi_7x28 multi_7x28_mod_1628(clk,rst,matrix_A[1628],matrix_B[28],mul_res1[1628]);
multi_7x28 multi_7x28_mod_1629(clk,rst,matrix_A[1629],matrix_B[29],mul_res1[1629]);
multi_7x28 multi_7x28_mod_1630(clk,rst,matrix_A[1630],matrix_B[30],mul_res1[1630]);
multi_7x28 multi_7x28_mod_1631(clk,rst,matrix_A[1631],matrix_B[31],mul_res1[1631]);
multi_7x28 multi_7x28_mod_1632(clk,rst,matrix_A[1632],matrix_B[32],mul_res1[1632]);
multi_7x28 multi_7x28_mod_1633(clk,rst,matrix_A[1633],matrix_B[33],mul_res1[1633]);
multi_7x28 multi_7x28_mod_1634(clk,rst,matrix_A[1634],matrix_B[34],mul_res1[1634]);
multi_7x28 multi_7x28_mod_1635(clk,rst,matrix_A[1635],matrix_B[35],mul_res1[1635]);
multi_7x28 multi_7x28_mod_1636(clk,rst,matrix_A[1636],matrix_B[36],mul_res1[1636]);
multi_7x28 multi_7x28_mod_1637(clk,rst,matrix_A[1637],matrix_B[37],mul_res1[1637]);
multi_7x28 multi_7x28_mod_1638(clk,rst,matrix_A[1638],matrix_B[38],mul_res1[1638]);
multi_7x28 multi_7x28_mod_1639(clk,rst,matrix_A[1639],matrix_B[39],mul_res1[1639]);
multi_7x28 multi_7x28_mod_1640(clk,rst,matrix_A[1640],matrix_B[40],mul_res1[1640]);
multi_7x28 multi_7x28_mod_1641(clk,rst,matrix_A[1641],matrix_B[41],mul_res1[1641]);
multi_7x28 multi_7x28_mod_1642(clk,rst,matrix_A[1642],matrix_B[42],mul_res1[1642]);
multi_7x28 multi_7x28_mod_1643(clk,rst,matrix_A[1643],matrix_B[43],mul_res1[1643]);
multi_7x28 multi_7x28_mod_1644(clk,rst,matrix_A[1644],matrix_B[44],mul_res1[1644]);
multi_7x28 multi_7x28_mod_1645(clk,rst,matrix_A[1645],matrix_B[45],mul_res1[1645]);
multi_7x28 multi_7x28_mod_1646(clk,rst,matrix_A[1646],matrix_B[46],mul_res1[1646]);
multi_7x28 multi_7x28_mod_1647(clk,rst,matrix_A[1647],matrix_B[47],mul_res1[1647]);
multi_7x28 multi_7x28_mod_1648(clk,rst,matrix_A[1648],matrix_B[48],mul_res1[1648]);
multi_7x28 multi_7x28_mod_1649(clk,rst,matrix_A[1649],matrix_B[49],mul_res1[1649]);
multi_7x28 multi_7x28_mod_1650(clk,rst,matrix_A[1650],matrix_B[50],mul_res1[1650]);
multi_7x28 multi_7x28_mod_1651(clk,rst,matrix_A[1651],matrix_B[51],mul_res1[1651]);
multi_7x28 multi_7x28_mod_1652(clk,rst,matrix_A[1652],matrix_B[52],mul_res1[1652]);
multi_7x28 multi_7x28_mod_1653(clk,rst,matrix_A[1653],matrix_B[53],mul_res1[1653]);
multi_7x28 multi_7x28_mod_1654(clk,rst,matrix_A[1654],matrix_B[54],mul_res1[1654]);
multi_7x28 multi_7x28_mod_1655(clk,rst,matrix_A[1655],matrix_B[55],mul_res1[1655]);
multi_7x28 multi_7x28_mod_1656(clk,rst,matrix_A[1656],matrix_B[56],mul_res1[1656]);
multi_7x28 multi_7x28_mod_1657(clk,rst,matrix_A[1657],matrix_B[57],mul_res1[1657]);
multi_7x28 multi_7x28_mod_1658(clk,rst,matrix_A[1658],matrix_B[58],mul_res1[1658]);
multi_7x28 multi_7x28_mod_1659(clk,rst,matrix_A[1659],matrix_B[59],mul_res1[1659]);
multi_7x28 multi_7x28_mod_1660(clk,rst,matrix_A[1660],matrix_B[60],mul_res1[1660]);
multi_7x28 multi_7x28_mod_1661(clk,rst,matrix_A[1661],matrix_B[61],mul_res1[1661]);
multi_7x28 multi_7x28_mod_1662(clk,rst,matrix_A[1662],matrix_B[62],mul_res1[1662]);
multi_7x28 multi_7x28_mod_1663(clk,rst,matrix_A[1663],matrix_B[63],mul_res1[1663]);
multi_7x28 multi_7x28_mod_1664(clk,rst,matrix_A[1664],matrix_B[64],mul_res1[1664]);
multi_7x28 multi_7x28_mod_1665(clk,rst,matrix_A[1665],matrix_B[65],mul_res1[1665]);
multi_7x28 multi_7x28_mod_1666(clk,rst,matrix_A[1666],matrix_B[66],mul_res1[1666]);
multi_7x28 multi_7x28_mod_1667(clk,rst,matrix_A[1667],matrix_B[67],mul_res1[1667]);
multi_7x28 multi_7x28_mod_1668(clk,rst,matrix_A[1668],matrix_B[68],mul_res1[1668]);
multi_7x28 multi_7x28_mod_1669(clk,rst,matrix_A[1669],matrix_B[69],mul_res1[1669]);
multi_7x28 multi_7x28_mod_1670(clk,rst,matrix_A[1670],matrix_B[70],mul_res1[1670]);
multi_7x28 multi_7x28_mod_1671(clk,rst,matrix_A[1671],matrix_B[71],mul_res1[1671]);
multi_7x28 multi_7x28_mod_1672(clk,rst,matrix_A[1672],matrix_B[72],mul_res1[1672]);
multi_7x28 multi_7x28_mod_1673(clk,rst,matrix_A[1673],matrix_B[73],mul_res1[1673]);
multi_7x28 multi_7x28_mod_1674(clk,rst,matrix_A[1674],matrix_B[74],mul_res1[1674]);
multi_7x28 multi_7x28_mod_1675(clk,rst,matrix_A[1675],matrix_B[75],mul_res1[1675]);
multi_7x28 multi_7x28_mod_1676(clk,rst,matrix_A[1676],matrix_B[76],mul_res1[1676]);
multi_7x28 multi_7x28_mod_1677(clk,rst,matrix_A[1677],matrix_B[77],mul_res1[1677]);
multi_7x28 multi_7x28_mod_1678(clk,rst,matrix_A[1678],matrix_B[78],mul_res1[1678]);
multi_7x28 multi_7x28_mod_1679(clk,rst,matrix_A[1679],matrix_B[79],mul_res1[1679]);
multi_7x28 multi_7x28_mod_1680(clk,rst,matrix_A[1680],matrix_B[80],mul_res1[1680]);
multi_7x28 multi_7x28_mod_1681(clk,rst,matrix_A[1681],matrix_B[81],mul_res1[1681]);
multi_7x28 multi_7x28_mod_1682(clk,rst,matrix_A[1682],matrix_B[82],mul_res1[1682]);
multi_7x28 multi_7x28_mod_1683(clk,rst,matrix_A[1683],matrix_B[83],mul_res1[1683]);
multi_7x28 multi_7x28_mod_1684(clk,rst,matrix_A[1684],matrix_B[84],mul_res1[1684]);
multi_7x28 multi_7x28_mod_1685(clk,rst,matrix_A[1685],matrix_B[85],mul_res1[1685]);
multi_7x28 multi_7x28_mod_1686(clk,rst,matrix_A[1686],matrix_B[86],mul_res1[1686]);
multi_7x28 multi_7x28_mod_1687(clk,rst,matrix_A[1687],matrix_B[87],mul_res1[1687]);
multi_7x28 multi_7x28_mod_1688(clk,rst,matrix_A[1688],matrix_B[88],mul_res1[1688]);
multi_7x28 multi_7x28_mod_1689(clk,rst,matrix_A[1689],matrix_B[89],mul_res1[1689]);
multi_7x28 multi_7x28_mod_1690(clk,rst,matrix_A[1690],matrix_B[90],mul_res1[1690]);
multi_7x28 multi_7x28_mod_1691(clk,rst,matrix_A[1691],matrix_B[91],mul_res1[1691]);
multi_7x28 multi_7x28_mod_1692(clk,rst,matrix_A[1692],matrix_B[92],mul_res1[1692]);
multi_7x28 multi_7x28_mod_1693(clk,rst,matrix_A[1693],matrix_B[93],mul_res1[1693]);
multi_7x28 multi_7x28_mod_1694(clk,rst,matrix_A[1694],matrix_B[94],mul_res1[1694]);
multi_7x28 multi_7x28_mod_1695(clk,rst,matrix_A[1695],matrix_B[95],mul_res1[1695]);
multi_7x28 multi_7x28_mod_1696(clk,rst,matrix_A[1696],matrix_B[96],mul_res1[1696]);
multi_7x28 multi_7x28_mod_1697(clk,rst,matrix_A[1697],matrix_B[97],mul_res1[1697]);
multi_7x28 multi_7x28_mod_1698(clk,rst,matrix_A[1698],matrix_B[98],mul_res1[1698]);
multi_7x28 multi_7x28_mod_1699(clk,rst,matrix_A[1699],matrix_B[99],mul_res1[1699]);
multi_7x28 multi_7x28_mod_1700(clk,rst,matrix_A[1700],matrix_B[100],mul_res1[1700]);
multi_7x28 multi_7x28_mod_1701(clk,rst,matrix_A[1701],matrix_B[101],mul_res1[1701]);
multi_7x28 multi_7x28_mod_1702(clk,rst,matrix_A[1702],matrix_B[102],mul_res1[1702]);
multi_7x28 multi_7x28_mod_1703(clk,rst,matrix_A[1703],matrix_B[103],mul_res1[1703]);
multi_7x28 multi_7x28_mod_1704(clk,rst,matrix_A[1704],matrix_B[104],mul_res1[1704]);
multi_7x28 multi_7x28_mod_1705(clk,rst,matrix_A[1705],matrix_B[105],mul_res1[1705]);
multi_7x28 multi_7x28_mod_1706(clk,rst,matrix_A[1706],matrix_B[106],mul_res1[1706]);
multi_7x28 multi_7x28_mod_1707(clk,rst,matrix_A[1707],matrix_B[107],mul_res1[1707]);
multi_7x28 multi_7x28_mod_1708(clk,rst,matrix_A[1708],matrix_B[108],mul_res1[1708]);
multi_7x28 multi_7x28_mod_1709(clk,rst,matrix_A[1709],matrix_B[109],mul_res1[1709]);
multi_7x28 multi_7x28_mod_1710(clk,rst,matrix_A[1710],matrix_B[110],mul_res1[1710]);
multi_7x28 multi_7x28_mod_1711(clk,rst,matrix_A[1711],matrix_B[111],mul_res1[1711]);
multi_7x28 multi_7x28_mod_1712(clk,rst,matrix_A[1712],matrix_B[112],mul_res1[1712]);
multi_7x28 multi_7x28_mod_1713(clk,rst,matrix_A[1713],matrix_B[113],mul_res1[1713]);
multi_7x28 multi_7x28_mod_1714(clk,rst,matrix_A[1714],matrix_B[114],mul_res1[1714]);
multi_7x28 multi_7x28_mod_1715(clk,rst,matrix_A[1715],matrix_B[115],mul_res1[1715]);
multi_7x28 multi_7x28_mod_1716(clk,rst,matrix_A[1716],matrix_B[116],mul_res1[1716]);
multi_7x28 multi_7x28_mod_1717(clk,rst,matrix_A[1717],matrix_B[117],mul_res1[1717]);
multi_7x28 multi_7x28_mod_1718(clk,rst,matrix_A[1718],matrix_B[118],mul_res1[1718]);
multi_7x28 multi_7x28_mod_1719(clk,rst,matrix_A[1719],matrix_B[119],mul_res1[1719]);
multi_7x28 multi_7x28_mod_1720(clk,rst,matrix_A[1720],matrix_B[120],mul_res1[1720]);
multi_7x28 multi_7x28_mod_1721(clk,rst,matrix_A[1721],matrix_B[121],mul_res1[1721]);
multi_7x28 multi_7x28_mod_1722(clk,rst,matrix_A[1722],matrix_B[122],mul_res1[1722]);
multi_7x28 multi_7x28_mod_1723(clk,rst,matrix_A[1723],matrix_B[123],mul_res1[1723]);
multi_7x28 multi_7x28_mod_1724(clk,rst,matrix_A[1724],matrix_B[124],mul_res1[1724]);
multi_7x28 multi_7x28_mod_1725(clk,rst,matrix_A[1725],matrix_B[125],mul_res1[1725]);
multi_7x28 multi_7x28_mod_1726(clk,rst,matrix_A[1726],matrix_B[126],mul_res1[1726]);
multi_7x28 multi_7x28_mod_1727(clk,rst,matrix_A[1727],matrix_B[127],mul_res1[1727]);
multi_7x28 multi_7x28_mod_1728(clk,rst,matrix_A[1728],matrix_B[128],mul_res1[1728]);
multi_7x28 multi_7x28_mod_1729(clk,rst,matrix_A[1729],matrix_B[129],mul_res1[1729]);
multi_7x28 multi_7x28_mod_1730(clk,rst,matrix_A[1730],matrix_B[130],mul_res1[1730]);
multi_7x28 multi_7x28_mod_1731(clk,rst,matrix_A[1731],matrix_B[131],mul_res1[1731]);
multi_7x28 multi_7x28_mod_1732(clk,rst,matrix_A[1732],matrix_B[132],mul_res1[1732]);
multi_7x28 multi_7x28_mod_1733(clk,rst,matrix_A[1733],matrix_B[133],mul_res1[1733]);
multi_7x28 multi_7x28_mod_1734(clk,rst,matrix_A[1734],matrix_B[134],mul_res1[1734]);
multi_7x28 multi_7x28_mod_1735(clk,rst,matrix_A[1735],matrix_B[135],mul_res1[1735]);
multi_7x28 multi_7x28_mod_1736(clk,rst,matrix_A[1736],matrix_B[136],mul_res1[1736]);
multi_7x28 multi_7x28_mod_1737(clk,rst,matrix_A[1737],matrix_B[137],mul_res1[1737]);
multi_7x28 multi_7x28_mod_1738(clk,rst,matrix_A[1738],matrix_B[138],mul_res1[1738]);
multi_7x28 multi_7x28_mod_1739(clk,rst,matrix_A[1739],matrix_B[139],mul_res1[1739]);
multi_7x28 multi_7x28_mod_1740(clk,rst,matrix_A[1740],matrix_B[140],mul_res1[1740]);
multi_7x28 multi_7x28_mod_1741(clk,rst,matrix_A[1741],matrix_B[141],mul_res1[1741]);
multi_7x28 multi_7x28_mod_1742(clk,rst,matrix_A[1742],matrix_B[142],mul_res1[1742]);
multi_7x28 multi_7x28_mod_1743(clk,rst,matrix_A[1743],matrix_B[143],mul_res1[1743]);
multi_7x28 multi_7x28_mod_1744(clk,rst,matrix_A[1744],matrix_B[144],mul_res1[1744]);
multi_7x28 multi_7x28_mod_1745(clk,rst,matrix_A[1745],matrix_B[145],mul_res1[1745]);
multi_7x28 multi_7x28_mod_1746(clk,rst,matrix_A[1746],matrix_B[146],mul_res1[1746]);
multi_7x28 multi_7x28_mod_1747(clk,rst,matrix_A[1747],matrix_B[147],mul_res1[1747]);
multi_7x28 multi_7x28_mod_1748(clk,rst,matrix_A[1748],matrix_B[148],mul_res1[1748]);
multi_7x28 multi_7x28_mod_1749(clk,rst,matrix_A[1749],matrix_B[149],mul_res1[1749]);
multi_7x28 multi_7x28_mod_1750(clk,rst,matrix_A[1750],matrix_B[150],mul_res1[1750]);
multi_7x28 multi_7x28_mod_1751(clk,rst,matrix_A[1751],matrix_B[151],mul_res1[1751]);
multi_7x28 multi_7x28_mod_1752(clk,rst,matrix_A[1752],matrix_B[152],mul_res1[1752]);
multi_7x28 multi_7x28_mod_1753(clk,rst,matrix_A[1753],matrix_B[153],mul_res1[1753]);
multi_7x28 multi_7x28_mod_1754(clk,rst,matrix_A[1754],matrix_B[154],mul_res1[1754]);
multi_7x28 multi_7x28_mod_1755(clk,rst,matrix_A[1755],matrix_B[155],mul_res1[1755]);
multi_7x28 multi_7x28_mod_1756(clk,rst,matrix_A[1756],matrix_B[156],mul_res1[1756]);
multi_7x28 multi_7x28_mod_1757(clk,rst,matrix_A[1757],matrix_B[157],mul_res1[1757]);
multi_7x28 multi_7x28_mod_1758(clk,rst,matrix_A[1758],matrix_B[158],mul_res1[1758]);
multi_7x28 multi_7x28_mod_1759(clk,rst,matrix_A[1759],matrix_B[159],mul_res1[1759]);
multi_7x28 multi_7x28_mod_1760(clk,rst,matrix_A[1760],matrix_B[160],mul_res1[1760]);
multi_7x28 multi_7x28_mod_1761(clk,rst,matrix_A[1761],matrix_B[161],mul_res1[1761]);
multi_7x28 multi_7x28_mod_1762(clk,rst,matrix_A[1762],matrix_B[162],mul_res1[1762]);
multi_7x28 multi_7x28_mod_1763(clk,rst,matrix_A[1763],matrix_B[163],mul_res1[1763]);
multi_7x28 multi_7x28_mod_1764(clk,rst,matrix_A[1764],matrix_B[164],mul_res1[1764]);
multi_7x28 multi_7x28_mod_1765(clk,rst,matrix_A[1765],matrix_B[165],mul_res1[1765]);
multi_7x28 multi_7x28_mod_1766(clk,rst,matrix_A[1766],matrix_B[166],mul_res1[1766]);
multi_7x28 multi_7x28_mod_1767(clk,rst,matrix_A[1767],matrix_B[167],mul_res1[1767]);
multi_7x28 multi_7x28_mod_1768(clk,rst,matrix_A[1768],matrix_B[168],mul_res1[1768]);
multi_7x28 multi_7x28_mod_1769(clk,rst,matrix_A[1769],matrix_B[169],mul_res1[1769]);
multi_7x28 multi_7x28_mod_1770(clk,rst,matrix_A[1770],matrix_B[170],mul_res1[1770]);
multi_7x28 multi_7x28_mod_1771(clk,rst,matrix_A[1771],matrix_B[171],mul_res1[1771]);
multi_7x28 multi_7x28_mod_1772(clk,rst,matrix_A[1772],matrix_B[172],mul_res1[1772]);
multi_7x28 multi_7x28_mod_1773(clk,rst,matrix_A[1773],matrix_B[173],mul_res1[1773]);
multi_7x28 multi_7x28_mod_1774(clk,rst,matrix_A[1774],matrix_B[174],mul_res1[1774]);
multi_7x28 multi_7x28_mod_1775(clk,rst,matrix_A[1775],matrix_B[175],mul_res1[1775]);
multi_7x28 multi_7x28_mod_1776(clk,rst,matrix_A[1776],matrix_B[176],mul_res1[1776]);
multi_7x28 multi_7x28_mod_1777(clk,rst,matrix_A[1777],matrix_B[177],mul_res1[1777]);
multi_7x28 multi_7x28_mod_1778(clk,rst,matrix_A[1778],matrix_B[178],mul_res1[1778]);
multi_7x28 multi_7x28_mod_1779(clk,rst,matrix_A[1779],matrix_B[179],mul_res1[1779]);
multi_7x28 multi_7x28_mod_1780(clk,rst,matrix_A[1780],matrix_B[180],mul_res1[1780]);
multi_7x28 multi_7x28_mod_1781(clk,rst,matrix_A[1781],matrix_B[181],mul_res1[1781]);
multi_7x28 multi_7x28_mod_1782(clk,rst,matrix_A[1782],matrix_B[182],mul_res1[1782]);
multi_7x28 multi_7x28_mod_1783(clk,rst,matrix_A[1783],matrix_B[183],mul_res1[1783]);
multi_7x28 multi_7x28_mod_1784(clk,rst,matrix_A[1784],matrix_B[184],mul_res1[1784]);
multi_7x28 multi_7x28_mod_1785(clk,rst,matrix_A[1785],matrix_B[185],mul_res1[1785]);
multi_7x28 multi_7x28_mod_1786(clk,rst,matrix_A[1786],matrix_B[186],mul_res1[1786]);
multi_7x28 multi_7x28_mod_1787(clk,rst,matrix_A[1787],matrix_B[187],mul_res1[1787]);
multi_7x28 multi_7x28_mod_1788(clk,rst,matrix_A[1788],matrix_B[188],mul_res1[1788]);
multi_7x28 multi_7x28_mod_1789(clk,rst,matrix_A[1789],matrix_B[189],mul_res1[1789]);
multi_7x28 multi_7x28_mod_1790(clk,rst,matrix_A[1790],matrix_B[190],mul_res1[1790]);
multi_7x28 multi_7x28_mod_1791(clk,rst,matrix_A[1791],matrix_B[191],mul_res1[1791]);
multi_7x28 multi_7x28_mod_1792(clk,rst,matrix_A[1792],matrix_B[192],mul_res1[1792]);
multi_7x28 multi_7x28_mod_1793(clk,rst,matrix_A[1793],matrix_B[193],mul_res1[1793]);
multi_7x28 multi_7x28_mod_1794(clk,rst,matrix_A[1794],matrix_B[194],mul_res1[1794]);
multi_7x28 multi_7x28_mod_1795(clk,rst,matrix_A[1795],matrix_B[195],mul_res1[1795]);
multi_7x28 multi_7x28_mod_1796(clk,rst,matrix_A[1796],matrix_B[196],mul_res1[1796]);
multi_7x28 multi_7x28_mod_1797(clk,rst,matrix_A[1797],matrix_B[197],mul_res1[1797]);
multi_7x28 multi_7x28_mod_1798(clk,rst,matrix_A[1798],matrix_B[198],mul_res1[1798]);
multi_7x28 multi_7x28_mod_1799(clk,rst,matrix_A[1799],matrix_B[199],mul_res1[1799]);
multi_7x28 multi_7x28_mod_1800(clk,rst,matrix_A[1800],matrix_B[0],mul_res1[1800]);
multi_7x28 multi_7x28_mod_1801(clk,rst,matrix_A[1801],matrix_B[1],mul_res1[1801]);
multi_7x28 multi_7x28_mod_1802(clk,rst,matrix_A[1802],matrix_B[2],mul_res1[1802]);
multi_7x28 multi_7x28_mod_1803(clk,rst,matrix_A[1803],matrix_B[3],mul_res1[1803]);
multi_7x28 multi_7x28_mod_1804(clk,rst,matrix_A[1804],matrix_B[4],mul_res1[1804]);
multi_7x28 multi_7x28_mod_1805(clk,rst,matrix_A[1805],matrix_B[5],mul_res1[1805]);
multi_7x28 multi_7x28_mod_1806(clk,rst,matrix_A[1806],matrix_B[6],mul_res1[1806]);
multi_7x28 multi_7x28_mod_1807(clk,rst,matrix_A[1807],matrix_B[7],mul_res1[1807]);
multi_7x28 multi_7x28_mod_1808(clk,rst,matrix_A[1808],matrix_B[8],mul_res1[1808]);
multi_7x28 multi_7x28_mod_1809(clk,rst,matrix_A[1809],matrix_B[9],mul_res1[1809]);
multi_7x28 multi_7x28_mod_1810(clk,rst,matrix_A[1810],matrix_B[10],mul_res1[1810]);
multi_7x28 multi_7x28_mod_1811(clk,rst,matrix_A[1811],matrix_B[11],mul_res1[1811]);
multi_7x28 multi_7x28_mod_1812(clk,rst,matrix_A[1812],matrix_B[12],mul_res1[1812]);
multi_7x28 multi_7x28_mod_1813(clk,rst,matrix_A[1813],matrix_B[13],mul_res1[1813]);
multi_7x28 multi_7x28_mod_1814(clk,rst,matrix_A[1814],matrix_B[14],mul_res1[1814]);
multi_7x28 multi_7x28_mod_1815(clk,rst,matrix_A[1815],matrix_B[15],mul_res1[1815]);
multi_7x28 multi_7x28_mod_1816(clk,rst,matrix_A[1816],matrix_B[16],mul_res1[1816]);
multi_7x28 multi_7x28_mod_1817(clk,rst,matrix_A[1817],matrix_B[17],mul_res1[1817]);
multi_7x28 multi_7x28_mod_1818(clk,rst,matrix_A[1818],matrix_B[18],mul_res1[1818]);
multi_7x28 multi_7x28_mod_1819(clk,rst,matrix_A[1819],matrix_B[19],mul_res1[1819]);
multi_7x28 multi_7x28_mod_1820(clk,rst,matrix_A[1820],matrix_B[20],mul_res1[1820]);
multi_7x28 multi_7x28_mod_1821(clk,rst,matrix_A[1821],matrix_B[21],mul_res1[1821]);
multi_7x28 multi_7x28_mod_1822(clk,rst,matrix_A[1822],matrix_B[22],mul_res1[1822]);
multi_7x28 multi_7x28_mod_1823(clk,rst,matrix_A[1823],matrix_B[23],mul_res1[1823]);
multi_7x28 multi_7x28_mod_1824(clk,rst,matrix_A[1824],matrix_B[24],mul_res1[1824]);
multi_7x28 multi_7x28_mod_1825(clk,rst,matrix_A[1825],matrix_B[25],mul_res1[1825]);
multi_7x28 multi_7x28_mod_1826(clk,rst,matrix_A[1826],matrix_B[26],mul_res1[1826]);
multi_7x28 multi_7x28_mod_1827(clk,rst,matrix_A[1827],matrix_B[27],mul_res1[1827]);
multi_7x28 multi_7x28_mod_1828(clk,rst,matrix_A[1828],matrix_B[28],mul_res1[1828]);
multi_7x28 multi_7x28_mod_1829(clk,rst,matrix_A[1829],matrix_B[29],mul_res1[1829]);
multi_7x28 multi_7x28_mod_1830(clk,rst,matrix_A[1830],matrix_B[30],mul_res1[1830]);
multi_7x28 multi_7x28_mod_1831(clk,rst,matrix_A[1831],matrix_B[31],mul_res1[1831]);
multi_7x28 multi_7x28_mod_1832(clk,rst,matrix_A[1832],matrix_B[32],mul_res1[1832]);
multi_7x28 multi_7x28_mod_1833(clk,rst,matrix_A[1833],matrix_B[33],mul_res1[1833]);
multi_7x28 multi_7x28_mod_1834(clk,rst,matrix_A[1834],matrix_B[34],mul_res1[1834]);
multi_7x28 multi_7x28_mod_1835(clk,rst,matrix_A[1835],matrix_B[35],mul_res1[1835]);
multi_7x28 multi_7x28_mod_1836(clk,rst,matrix_A[1836],matrix_B[36],mul_res1[1836]);
multi_7x28 multi_7x28_mod_1837(clk,rst,matrix_A[1837],matrix_B[37],mul_res1[1837]);
multi_7x28 multi_7x28_mod_1838(clk,rst,matrix_A[1838],matrix_B[38],mul_res1[1838]);
multi_7x28 multi_7x28_mod_1839(clk,rst,matrix_A[1839],matrix_B[39],mul_res1[1839]);
multi_7x28 multi_7x28_mod_1840(clk,rst,matrix_A[1840],matrix_B[40],mul_res1[1840]);
multi_7x28 multi_7x28_mod_1841(clk,rst,matrix_A[1841],matrix_B[41],mul_res1[1841]);
multi_7x28 multi_7x28_mod_1842(clk,rst,matrix_A[1842],matrix_B[42],mul_res1[1842]);
multi_7x28 multi_7x28_mod_1843(clk,rst,matrix_A[1843],matrix_B[43],mul_res1[1843]);
multi_7x28 multi_7x28_mod_1844(clk,rst,matrix_A[1844],matrix_B[44],mul_res1[1844]);
multi_7x28 multi_7x28_mod_1845(clk,rst,matrix_A[1845],matrix_B[45],mul_res1[1845]);
multi_7x28 multi_7x28_mod_1846(clk,rst,matrix_A[1846],matrix_B[46],mul_res1[1846]);
multi_7x28 multi_7x28_mod_1847(clk,rst,matrix_A[1847],matrix_B[47],mul_res1[1847]);
multi_7x28 multi_7x28_mod_1848(clk,rst,matrix_A[1848],matrix_B[48],mul_res1[1848]);
multi_7x28 multi_7x28_mod_1849(clk,rst,matrix_A[1849],matrix_B[49],mul_res1[1849]);
multi_7x28 multi_7x28_mod_1850(clk,rst,matrix_A[1850],matrix_B[50],mul_res1[1850]);
multi_7x28 multi_7x28_mod_1851(clk,rst,matrix_A[1851],matrix_B[51],mul_res1[1851]);
multi_7x28 multi_7x28_mod_1852(clk,rst,matrix_A[1852],matrix_B[52],mul_res1[1852]);
multi_7x28 multi_7x28_mod_1853(clk,rst,matrix_A[1853],matrix_B[53],mul_res1[1853]);
multi_7x28 multi_7x28_mod_1854(clk,rst,matrix_A[1854],matrix_B[54],mul_res1[1854]);
multi_7x28 multi_7x28_mod_1855(clk,rst,matrix_A[1855],matrix_B[55],mul_res1[1855]);
multi_7x28 multi_7x28_mod_1856(clk,rst,matrix_A[1856],matrix_B[56],mul_res1[1856]);
multi_7x28 multi_7x28_mod_1857(clk,rst,matrix_A[1857],matrix_B[57],mul_res1[1857]);
multi_7x28 multi_7x28_mod_1858(clk,rst,matrix_A[1858],matrix_B[58],mul_res1[1858]);
multi_7x28 multi_7x28_mod_1859(clk,rst,matrix_A[1859],matrix_B[59],mul_res1[1859]);
multi_7x28 multi_7x28_mod_1860(clk,rst,matrix_A[1860],matrix_B[60],mul_res1[1860]);
multi_7x28 multi_7x28_mod_1861(clk,rst,matrix_A[1861],matrix_B[61],mul_res1[1861]);
multi_7x28 multi_7x28_mod_1862(clk,rst,matrix_A[1862],matrix_B[62],mul_res1[1862]);
multi_7x28 multi_7x28_mod_1863(clk,rst,matrix_A[1863],matrix_B[63],mul_res1[1863]);
multi_7x28 multi_7x28_mod_1864(clk,rst,matrix_A[1864],matrix_B[64],mul_res1[1864]);
multi_7x28 multi_7x28_mod_1865(clk,rst,matrix_A[1865],matrix_B[65],mul_res1[1865]);
multi_7x28 multi_7x28_mod_1866(clk,rst,matrix_A[1866],matrix_B[66],mul_res1[1866]);
multi_7x28 multi_7x28_mod_1867(clk,rst,matrix_A[1867],matrix_B[67],mul_res1[1867]);
multi_7x28 multi_7x28_mod_1868(clk,rst,matrix_A[1868],matrix_B[68],mul_res1[1868]);
multi_7x28 multi_7x28_mod_1869(clk,rst,matrix_A[1869],matrix_B[69],mul_res1[1869]);
multi_7x28 multi_7x28_mod_1870(clk,rst,matrix_A[1870],matrix_B[70],mul_res1[1870]);
multi_7x28 multi_7x28_mod_1871(clk,rst,matrix_A[1871],matrix_B[71],mul_res1[1871]);
multi_7x28 multi_7x28_mod_1872(clk,rst,matrix_A[1872],matrix_B[72],mul_res1[1872]);
multi_7x28 multi_7x28_mod_1873(clk,rst,matrix_A[1873],matrix_B[73],mul_res1[1873]);
multi_7x28 multi_7x28_mod_1874(clk,rst,matrix_A[1874],matrix_B[74],mul_res1[1874]);
multi_7x28 multi_7x28_mod_1875(clk,rst,matrix_A[1875],matrix_B[75],mul_res1[1875]);
multi_7x28 multi_7x28_mod_1876(clk,rst,matrix_A[1876],matrix_B[76],mul_res1[1876]);
multi_7x28 multi_7x28_mod_1877(clk,rst,matrix_A[1877],matrix_B[77],mul_res1[1877]);
multi_7x28 multi_7x28_mod_1878(clk,rst,matrix_A[1878],matrix_B[78],mul_res1[1878]);
multi_7x28 multi_7x28_mod_1879(clk,rst,matrix_A[1879],matrix_B[79],mul_res1[1879]);
multi_7x28 multi_7x28_mod_1880(clk,rst,matrix_A[1880],matrix_B[80],mul_res1[1880]);
multi_7x28 multi_7x28_mod_1881(clk,rst,matrix_A[1881],matrix_B[81],mul_res1[1881]);
multi_7x28 multi_7x28_mod_1882(clk,rst,matrix_A[1882],matrix_B[82],mul_res1[1882]);
multi_7x28 multi_7x28_mod_1883(clk,rst,matrix_A[1883],matrix_B[83],mul_res1[1883]);
multi_7x28 multi_7x28_mod_1884(clk,rst,matrix_A[1884],matrix_B[84],mul_res1[1884]);
multi_7x28 multi_7x28_mod_1885(clk,rst,matrix_A[1885],matrix_B[85],mul_res1[1885]);
multi_7x28 multi_7x28_mod_1886(clk,rst,matrix_A[1886],matrix_B[86],mul_res1[1886]);
multi_7x28 multi_7x28_mod_1887(clk,rst,matrix_A[1887],matrix_B[87],mul_res1[1887]);
multi_7x28 multi_7x28_mod_1888(clk,rst,matrix_A[1888],matrix_B[88],mul_res1[1888]);
multi_7x28 multi_7x28_mod_1889(clk,rst,matrix_A[1889],matrix_B[89],mul_res1[1889]);
multi_7x28 multi_7x28_mod_1890(clk,rst,matrix_A[1890],matrix_B[90],mul_res1[1890]);
multi_7x28 multi_7x28_mod_1891(clk,rst,matrix_A[1891],matrix_B[91],mul_res1[1891]);
multi_7x28 multi_7x28_mod_1892(clk,rst,matrix_A[1892],matrix_B[92],mul_res1[1892]);
multi_7x28 multi_7x28_mod_1893(clk,rst,matrix_A[1893],matrix_B[93],mul_res1[1893]);
multi_7x28 multi_7x28_mod_1894(clk,rst,matrix_A[1894],matrix_B[94],mul_res1[1894]);
multi_7x28 multi_7x28_mod_1895(clk,rst,matrix_A[1895],matrix_B[95],mul_res1[1895]);
multi_7x28 multi_7x28_mod_1896(clk,rst,matrix_A[1896],matrix_B[96],mul_res1[1896]);
multi_7x28 multi_7x28_mod_1897(clk,rst,matrix_A[1897],matrix_B[97],mul_res1[1897]);
multi_7x28 multi_7x28_mod_1898(clk,rst,matrix_A[1898],matrix_B[98],mul_res1[1898]);
multi_7x28 multi_7x28_mod_1899(clk,rst,matrix_A[1899],matrix_B[99],mul_res1[1899]);
multi_7x28 multi_7x28_mod_1900(clk,rst,matrix_A[1900],matrix_B[100],mul_res1[1900]);
multi_7x28 multi_7x28_mod_1901(clk,rst,matrix_A[1901],matrix_B[101],mul_res1[1901]);
multi_7x28 multi_7x28_mod_1902(clk,rst,matrix_A[1902],matrix_B[102],mul_res1[1902]);
multi_7x28 multi_7x28_mod_1903(clk,rst,matrix_A[1903],matrix_B[103],mul_res1[1903]);
multi_7x28 multi_7x28_mod_1904(clk,rst,matrix_A[1904],matrix_B[104],mul_res1[1904]);
multi_7x28 multi_7x28_mod_1905(clk,rst,matrix_A[1905],matrix_B[105],mul_res1[1905]);
multi_7x28 multi_7x28_mod_1906(clk,rst,matrix_A[1906],matrix_B[106],mul_res1[1906]);
multi_7x28 multi_7x28_mod_1907(clk,rst,matrix_A[1907],matrix_B[107],mul_res1[1907]);
multi_7x28 multi_7x28_mod_1908(clk,rst,matrix_A[1908],matrix_B[108],mul_res1[1908]);
multi_7x28 multi_7x28_mod_1909(clk,rst,matrix_A[1909],matrix_B[109],mul_res1[1909]);
multi_7x28 multi_7x28_mod_1910(clk,rst,matrix_A[1910],matrix_B[110],mul_res1[1910]);
multi_7x28 multi_7x28_mod_1911(clk,rst,matrix_A[1911],matrix_B[111],mul_res1[1911]);
multi_7x28 multi_7x28_mod_1912(clk,rst,matrix_A[1912],matrix_B[112],mul_res1[1912]);
multi_7x28 multi_7x28_mod_1913(clk,rst,matrix_A[1913],matrix_B[113],mul_res1[1913]);
multi_7x28 multi_7x28_mod_1914(clk,rst,matrix_A[1914],matrix_B[114],mul_res1[1914]);
multi_7x28 multi_7x28_mod_1915(clk,rst,matrix_A[1915],matrix_B[115],mul_res1[1915]);
multi_7x28 multi_7x28_mod_1916(clk,rst,matrix_A[1916],matrix_B[116],mul_res1[1916]);
multi_7x28 multi_7x28_mod_1917(clk,rst,matrix_A[1917],matrix_B[117],mul_res1[1917]);
multi_7x28 multi_7x28_mod_1918(clk,rst,matrix_A[1918],matrix_B[118],mul_res1[1918]);
multi_7x28 multi_7x28_mod_1919(clk,rst,matrix_A[1919],matrix_B[119],mul_res1[1919]);
multi_7x28 multi_7x28_mod_1920(clk,rst,matrix_A[1920],matrix_B[120],mul_res1[1920]);
multi_7x28 multi_7x28_mod_1921(clk,rst,matrix_A[1921],matrix_B[121],mul_res1[1921]);
multi_7x28 multi_7x28_mod_1922(clk,rst,matrix_A[1922],matrix_B[122],mul_res1[1922]);
multi_7x28 multi_7x28_mod_1923(clk,rst,matrix_A[1923],matrix_B[123],mul_res1[1923]);
multi_7x28 multi_7x28_mod_1924(clk,rst,matrix_A[1924],matrix_B[124],mul_res1[1924]);
multi_7x28 multi_7x28_mod_1925(clk,rst,matrix_A[1925],matrix_B[125],mul_res1[1925]);
multi_7x28 multi_7x28_mod_1926(clk,rst,matrix_A[1926],matrix_B[126],mul_res1[1926]);
multi_7x28 multi_7x28_mod_1927(clk,rst,matrix_A[1927],matrix_B[127],mul_res1[1927]);
multi_7x28 multi_7x28_mod_1928(clk,rst,matrix_A[1928],matrix_B[128],mul_res1[1928]);
multi_7x28 multi_7x28_mod_1929(clk,rst,matrix_A[1929],matrix_B[129],mul_res1[1929]);
multi_7x28 multi_7x28_mod_1930(clk,rst,matrix_A[1930],matrix_B[130],mul_res1[1930]);
multi_7x28 multi_7x28_mod_1931(clk,rst,matrix_A[1931],matrix_B[131],mul_res1[1931]);
multi_7x28 multi_7x28_mod_1932(clk,rst,matrix_A[1932],matrix_B[132],mul_res1[1932]);
multi_7x28 multi_7x28_mod_1933(clk,rst,matrix_A[1933],matrix_B[133],mul_res1[1933]);
multi_7x28 multi_7x28_mod_1934(clk,rst,matrix_A[1934],matrix_B[134],mul_res1[1934]);
multi_7x28 multi_7x28_mod_1935(clk,rst,matrix_A[1935],matrix_B[135],mul_res1[1935]);
multi_7x28 multi_7x28_mod_1936(clk,rst,matrix_A[1936],matrix_B[136],mul_res1[1936]);
multi_7x28 multi_7x28_mod_1937(clk,rst,matrix_A[1937],matrix_B[137],mul_res1[1937]);
multi_7x28 multi_7x28_mod_1938(clk,rst,matrix_A[1938],matrix_B[138],mul_res1[1938]);
multi_7x28 multi_7x28_mod_1939(clk,rst,matrix_A[1939],matrix_B[139],mul_res1[1939]);
multi_7x28 multi_7x28_mod_1940(clk,rst,matrix_A[1940],matrix_B[140],mul_res1[1940]);
multi_7x28 multi_7x28_mod_1941(clk,rst,matrix_A[1941],matrix_B[141],mul_res1[1941]);
multi_7x28 multi_7x28_mod_1942(clk,rst,matrix_A[1942],matrix_B[142],mul_res1[1942]);
multi_7x28 multi_7x28_mod_1943(clk,rst,matrix_A[1943],matrix_B[143],mul_res1[1943]);
multi_7x28 multi_7x28_mod_1944(clk,rst,matrix_A[1944],matrix_B[144],mul_res1[1944]);
multi_7x28 multi_7x28_mod_1945(clk,rst,matrix_A[1945],matrix_B[145],mul_res1[1945]);
multi_7x28 multi_7x28_mod_1946(clk,rst,matrix_A[1946],matrix_B[146],mul_res1[1946]);
multi_7x28 multi_7x28_mod_1947(clk,rst,matrix_A[1947],matrix_B[147],mul_res1[1947]);
multi_7x28 multi_7x28_mod_1948(clk,rst,matrix_A[1948],matrix_B[148],mul_res1[1948]);
multi_7x28 multi_7x28_mod_1949(clk,rst,matrix_A[1949],matrix_B[149],mul_res1[1949]);
multi_7x28 multi_7x28_mod_1950(clk,rst,matrix_A[1950],matrix_B[150],mul_res1[1950]);
multi_7x28 multi_7x28_mod_1951(clk,rst,matrix_A[1951],matrix_B[151],mul_res1[1951]);
multi_7x28 multi_7x28_mod_1952(clk,rst,matrix_A[1952],matrix_B[152],mul_res1[1952]);
multi_7x28 multi_7x28_mod_1953(clk,rst,matrix_A[1953],matrix_B[153],mul_res1[1953]);
multi_7x28 multi_7x28_mod_1954(clk,rst,matrix_A[1954],matrix_B[154],mul_res1[1954]);
multi_7x28 multi_7x28_mod_1955(clk,rst,matrix_A[1955],matrix_B[155],mul_res1[1955]);
multi_7x28 multi_7x28_mod_1956(clk,rst,matrix_A[1956],matrix_B[156],mul_res1[1956]);
multi_7x28 multi_7x28_mod_1957(clk,rst,matrix_A[1957],matrix_B[157],mul_res1[1957]);
multi_7x28 multi_7x28_mod_1958(clk,rst,matrix_A[1958],matrix_B[158],mul_res1[1958]);
multi_7x28 multi_7x28_mod_1959(clk,rst,matrix_A[1959],matrix_B[159],mul_res1[1959]);
multi_7x28 multi_7x28_mod_1960(clk,rst,matrix_A[1960],matrix_B[160],mul_res1[1960]);
multi_7x28 multi_7x28_mod_1961(clk,rst,matrix_A[1961],matrix_B[161],mul_res1[1961]);
multi_7x28 multi_7x28_mod_1962(clk,rst,matrix_A[1962],matrix_B[162],mul_res1[1962]);
multi_7x28 multi_7x28_mod_1963(clk,rst,matrix_A[1963],matrix_B[163],mul_res1[1963]);
multi_7x28 multi_7x28_mod_1964(clk,rst,matrix_A[1964],matrix_B[164],mul_res1[1964]);
multi_7x28 multi_7x28_mod_1965(clk,rst,matrix_A[1965],matrix_B[165],mul_res1[1965]);
multi_7x28 multi_7x28_mod_1966(clk,rst,matrix_A[1966],matrix_B[166],mul_res1[1966]);
multi_7x28 multi_7x28_mod_1967(clk,rst,matrix_A[1967],matrix_B[167],mul_res1[1967]);
multi_7x28 multi_7x28_mod_1968(clk,rst,matrix_A[1968],matrix_B[168],mul_res1[1968]);
multi_7x28 multi_7x28_mod_1969(clk,rst,matrix_A[1969],matrix_B[169],mul_res1[1969]);
multi_7x28 multi_7x28_mod_1970(clk,rst,matrix_A[1970],matrix_B[170],mul_res1[1970]);
multi_7x28 multi_7x28_mod_1971(clk,rst,matrix_A[1971],matrix_B[171],mul_res1[1971]);
multi_7x28 multi_7x28_mod_1972(clk,rst,matrix_A[1972],matrix_B[172],mul_res1[1972]);
multi_7x28 multi_7x28_mod_1973(clk,rst,matrix_A[1973],matrix_B[173],mul_res1[1973]);
multi_7x28 multi_7x28_mod_1974(clk,rst,matrix_A[1974],matrix_B[174],mul_res1[1974]);
multi_7x28 multi_7x28_mod_1975(clk,rst,matrix_A[1975],matrix_B[175],mul_res1[1975]);
multi_7x28 multi_7x28_mod_1976(clk,rst,matrix_A[1976],matrix_B[176],mul_res1[1976]);
multi_7x28 multi_7x28_mod_1977(clk,rst,matrix_A[1977],matrix_B[177],mul_res1[1977]);
multi_7x28 multi_7x28_mod_1978(clk,rst,matrix_A[1978],matrix_B[178],mul_res1[1978]);
multi_7x28 multi_7x28_mod_1979(clk,rst,matrix_A[1979],matrix_B[179],mul_res1[1979]);
multi_7x28 multi_7x28_mod_1980(clk,rst,matrix_A[1980],matrix_B[180],mul_res1[1980]);
multi_7x28 multi_7x28_mod_1981(clk,rst,matrix_A[1981],matrix_B[181],mul_res1[1981]);
multi_7x28 multi_7x28_mod_1982(clk,rst,matrix_A[1982],matrix_B[182],mul_res1[1982]);
multi_7x28 multi_7x28_mod_1983(clk,rst,matrix_A[1983],matrix_B[183],mul_res1[1983]);
multi_7x28 multi_7x28_mod_1984(clk,rst,matrix_A[1984],matrix_B[184],mul_res1[1984]);
multi_7x28 multi_7x28_mod_1985(clk,rst,matrix_A[1985],matrix_B[185],mul_res1[1985]);
multi_7x28 multi_7x28_mod_1986(clk,rst,matrix_A[1986],matrix_B[186],mul_res1[1986]);
multi_7x28 multi_7x28_mod_1987(clk,rst,matrix_A[1987],matrix_B[187],mul_res1[1987]);
multi_7x28 multi_7x28_mod_1988(clk,rst,matrix_A[1988],matrix_B[188],mul_res1[1988]);
multi_7x28 multi_7x28_mod_1989(clk,rst,matrix_A[1989],matrix_B[189],mul_res1[1989]);
multi_7x28 multi_7x28_mod_1990(clk,rst,matrix_A[1990],matrix_B[190],mul_res1[1990]);
multi_7x28 multi_7x28_mod_1991(clk,rst,matrix_A[1991],matrix_B[191],mul_res1[1991]);
multi_7x28 multi_7x28_mod_1992(clk,rst,matrix_A[1992],matrix_B[192],mul_res1[1992]);
multi_7x28 multi_7x28_mod_1993(clk,rst,matrix_A[1993],matrix_B[193],mul_res1[1993]);
multi_7x28 multi_7x28_mod_1994(clk,rst,matrix_A[1994],matrix_B[194],mul_res1[1994]);
multi_7x28 multi_7x28_mod_1995(clk,rst,matrix_A[1995],matrix_B[195],mul_res1[1995]);
multi_7x28 multi_7x28_mod_1996(clk,rst,matrix_A[1996],matrix_B[196],mul_res1[1996]);
multi_7x28 multi_7x28_mod_1997(clk,rst,matrix_A[1997],matrix_B[197],mul_res1[1997]);
multi_7x28 multi_7x28_mod_1998(clk,rst,matrix_A[1998],matrix_B[198],mul_res1[1998]);
multi_7x28 multi_7x28_mod_1999(clk,rst,matrix_A[1999],matrix_B[199],mul_res1[1999]);
multi_7x28 multi_7x28_mod_2000(clk,rst,matrix_A[2000],matrix_B[0],mul_res1[2000]);
multi_7x28 multi_7x28_mod_2001(clk,rst,matrix_A[2001],matrix_B[1],mul_res1[2001]);
multi_7x28 multi_7x28_mod_2002(clk,rst,matrix_A[2002],matrix_B[2],mul_res1[2002]);
multi_7x28 multi_7x28_mod_2003(clk,rst,matrix_A[2003],matrix_B[3],mul_res1[2003]);
multi_7x28 multi_7x28_mod_2004(clk,rst,matrix_A[2004],matrix_B[4],mul_res1[2004]);
multi_7x28 multi_7x28_mod_2005(clk,rst,matrix_A[2005],matrix_B[5],mul_res1[2005]);
multi_7x28 multi_7x28_mod_2006(clk,rst,matrix_A[2006],matrix_B[6],mul_res1[2006]);
multi_7x28 multi_7x28_mod_2007(clk,rst,matrix_A[2007],matrix_B[7],mul_res1[2007]);
multi_7x28 multi_7x28_mod_2008(clk,rst,matrix_A[2008],matrix_B[8],mul_res1[2008]);
multi_7x28 multi_7x28_mod_2009(clk,rst,matrix_A[2009],matrix_B[9],mul_res1[2009]);
multi_7x28 multi_7x28_mod_2010(clk,rst,matrix_A[2010],matrix_B[10],mul_res1[2010]);
multi_7x28 multi_7x28_mod_2011(clk,rst,matrix_A[2011],matrix_B[11],mul_res1[2011]);
multi_7x28 multi_7x28_mod_2012(clk,rst,matrix_A[2012],matrix_B[12],mul_res1[2012]);
multi_7x28 multi_7x28_mod_2013(clk,rst,matrix_A[2013],matrix_B[13],mul_res1[2013]);
multi_7x28 multi_7x28_mod_2014(clk,rst,matrix_A[2014],matrix_B[14],mul_res1[2014]);
multi_7x28 multi_7x28_mod_2015(clk,rst,matrix_A[2015],matrix_B[15],mul_res1[2015]);
multi_7x28 multi_7x28_mod_2016(clk,rst,matrix_A[2016],matrix_B[16],mul_res1[2016]);
multi_7x28 multi_7x28_mod_2017(clk,rst,matrix_A[2017],matrix_B[17],mul_res1[2017]);
multi_7x28 multi_7x28_mod_2018(clk,rst,matrix_A[2018],matrix_B[18],mul_res1[2018]);
multi_7x28 multi_7x28_mod_2019(clk,rst,matrix_A[2019],matrix_B[19],mul_res1[2019]);
multi_7x28 multi_7x28_mod_2020(clk,rst,matrix_A[2020],matrix_B[20],mul_res1[2020]);
multi_7x28 multi_7x28_mod_2021(clk,rst,matrix_A[2021],matrix_B[21],mul_res1[2021]);
multi_7x28 multi_7x28_mod_2022(clk,rst,matrix_A[2022],matrix_B[22],mul_res1[2022]);
multi_7x28 multi_7x28_mod_2023(clk,rst,matrix_A[2023],matrix_B[23],mul_res1[2023]);
multi_7x28 multi_7x28_mod_2024(clk,rst,matrix_A[2024],matrix_B[24],mul_res1[2024]);
multi_7x28 multi_7x28_mod_2025(clk,rst,matrix_A[2025],matrix_B[25],mul_res1[2025]);
multi_7x28 multi_7x28_mod_2026(clk,rst,matrix_A[2026],matrix_B[26],mul_res1[2026]);
multi_7x28 multi_7x28_mod_2027(clk,rst,matrix_A[2027],matrix_B[27],mul_res1[2027]);
multi_7x28 multi_7x28_mod_2028(clk,rst,matrix_A[2028],matrix_B[28],mul_res1[2028]);
multi_7x28 multi_7x28_mod_2029(clk,rst,matrix_A[2029],matrix_B[29],mul_res1[2029]);
multi_7x28 multi_7x28_mod_2030(clk,rst,matrix_A[2030],matrix_B[30],mul_res1[2030]);
multi_7x28 multi_7x28_mod_2031(clk,rst,matrix_A[2031],matrix_B[31],mul_res1[2031]);
multi_7x28 multi_7x28_mod_2032(clk,rst,matrix_A[2032],matrix_B[32],mul_res1[2032]);
multi_7x28 multi_7x28_mod_2033(clk,rst,matrix_A[2033],matrix_B[33],mul_res1[2033]);
multi_7x28 multi_7x28_mod_2034(clk,rst,matrix_A[2034],matrix_B[34],mul_res1[2034]);
multi_7x28 multi_7x28_mod_2035(clk,rst,matrix_A[2035],matrix_B[35],mul_res1[2035]);
multi_7x28 multi_7x28_mod_2036(clk,rst,matrix_A[2036],matrix_B[36],mul_res1[2036]);
multi_7x28 multi_7x28_mod_2037(clk,rst,matrix_A[2037],matrix_B[37],mul_res1[2037]);
multi_7x28 multi_7x28_mod_2038(clk,rst,matrix_A[2038],matrix_B[38],mul_res1[2038]);
multi_7x28 multi_7x28_mod_2039(clk,rst,matrix_A[2039],matrix_B[39],mul_res1[2039]);
multi_7x28 multi_7x28_mod_2040(clk,rst,matrix_A[2040],matrix_B[40],mul_res1[2040]);
multi_7x28 multi_7x28_mod_2041(clk,rst,matrix_A[2041],matrix_B[41],mul_res1[2041]);
multi_7x28 multi_7x28_mod_2042(clk,rst,matrix_A[2042],matrix_B[42],mul_res1[2042]);
multi_7x28 multi_7x28_mod_2043(clk,rst,matrix_A[2043],matrix_B[43],mul_res1[2043]);
multi_7x28 multi_7x28_mod_2044(clk,rst,matrix_A[2044],matrix_B[44],mul_res1[2044]);
multi_7x28 multi_7x28_mod_2045(clk,rst,matrix_A[2045],matrix_B[45],mul_res1[2045]);
multi_7x28 multi_7x28_mod_2046(clk,rst,matrix_A[2046],matrix_B[46],mul_res1[2046]);
multi_7x28 multi_7x28_mod_2047(clk,rst,matrix_A[2047],matrix_B[47],mul_res1[2047]);
multi_7x28 multi_7x28_mod_2048(clk,rst,matrix_A[2048],matrix_B[48],mul_res1[2048]);
multi_7x28 multi_7x28_mod_2049(clk,rst,matrix_A[2049],matrix_B[49],mul_res1[2049]);
multi_7x28 multi_7x28_mod_2050(clk,rst,matrix_A[2050],matrix_B[50],mul_res1[2050]);
multi_7x28 multi_7x28_mod_2051(clk,rst,matrix_A[2051],matrix_B[51],mul_res1[2051]);
multi_7x28 multi_7x28_mod_2052(clk,rst,matrix_A[2052],matrix_B[52],mul_res1[2052]);
multi_7x28 multi_7x28_mod_2053(clk,rst,matrix_A[2053],matrix_B[53],mul_res1[2053]);
multi_7x28 multi_7x28_mod_2054(clk,rst,matrix_A[2054],matrix_B[54],mul_res1[2054]);
multi_7x28 multi_7x28_mod_2055(clk,rst,matrix_A[2055],matrix_B[55],mul_res1[2055]);
multi_7x28 multi_7x28_mod_2056(clk,rst,matrix_A[2056],matrix_B[56],mul_res1[2056]);
multi_7x28 multi_7x28_mod_2057(clk,rst,matrix_A[2057],matrix_B[57],mul_res1[2057]);
multi_7x28 multi_7x28_mod_2058(clk,rst,matrix_A[2058],matrix_B[58],mul_res1[2058]);
multi_7x28 multi_7x28_mod_2059(clk,rst,matrix_A[2059],matrix_B[59],mul_res1[2059]);
multi_7x28 multi_7x28_mod_2060(clk,rst,matrix_A[2060],matrix_B[60],mul_res1[2060]);
multi_7x28 multi_7x28_mod_2061(clk,rst,matrix_A[2061],matrix_B[61],mul_res1[2061]);
multi_7x28 multi_7x28_mod_2062(clk,rst,matrix_A[2062],matrix_B[62],mul_res1[2062]);
multi_7x28 multi_7x28_mod_2063(clk,rst,matrix_A[2063],matrix_B[63],mul_res1[2063]);
multi_7x28 multi_7x28_mod_2064(clk,rst,matrix_A[2064],matrix_B[64],mul_res1[2064]);
multi_7x28 multi_7x28_mod_2065(clk,rst,matrix_A[2065],matrix_B[65],mul_res1[2065]);
multi_7x28 multi_7x28_mod_2066(clk,rst,matrix_A[2066],matrix_B[66],mul_res1[2066]);
multi_7x28 multi_7x28_mod_2067(clk,rst,matrix_A[2067],matrix_B[67],mul_res1[2067]);
multi_7x28 multi_7x28_mod_2068(clk,rst,matrix_A[2068],matrix_B[68],mul_res1[2068]);
multi_7x28 multi_7x28_mod_2069(clk,rst,matrix_A[2069],matrix_B[69],mul_res1[2069]);
multi_7x28 multi_7x28_mod_2070(clk,rst,matrix_A[2070],matrix_B[70],mul_res1[2070]);
multi_7x28 multi_7x28_mod_2071(clk,rst,matrix_A[2071],matrix_B[71],mul_res1[2071]);
multi_7x28 multi_7x28_mod_2072(clk,rst,matrix_A[2072],matrix_B[72],mul_res1[2072]);
multi_7x28 multi_7x28_mod_2073(clk,rst,matrix_A[2073],matrix_B[73],mul_res1[2073]);
multi_7x28 multi_7x28_mod_2074(clk,rst,matrix_A[2074],matrix_B[74],mul_res1[2074]);
multi_7x28 multi_7x28_mod_2075(clk,rst,matrix_A[2075],matrix_B[75],mul_res1[2075]);
multi_7x28 multi_7x28_mod_2076(clk,rst,matrix_A[2076],matrix_B[76],mul_res1[2076]);
multi_7x28 multi_7x28_mod_2077(clk,rst,matrix_A[2077],matrix_B[77],mul_res1[2077]);
multi_7x28 multi_7x28_mod_2078(clk,rst,matrix_A[2078],matrix_B[78],mul_res1[2078]);
multi_7x28 multi_7x28_mod_2079(clk,rst,matrix_A[2079],matrix_B[79],mul_res1[2079]);
multi_7x28 multi_7x28_mod_2080(clk,rst,matrix_A[2080],matrix_B[80],mul_res1[2080]);
multi_7x28 multi_7x28_mod_2081(clk,rst,matrix_A[2081],matrix_B[81],mul_res1[2081]);
multi_7x28 multi_7x28_mod_2082(clk,rst,matrix_A[2082],matrix_B[82],mul_res1[2082]);
multi_7x28 multi_7x28_mod_2083(clk,rst,matrix_A[2083],matrix_B[83],mul_res1[2083]);
multi_7x28 multi_7x28_mod_2084(clk,rst,matrix_A[2084],matrix_B[84],mul_res1[2084]);
multi_7x28 multi_7x28_mod_2085(clk,rst,matrix_A[2085],matrix_B[85],mul_res1[2085]);
multi_7x28 multi_7x28_mod_2086(clk,rst,matrix_A[2086],matrix_B[86],mul_res1[2086]);
multi_7x28 multi_7x28_mod_2087(clk,rst,matrix_A[2087],matrix_B[87],mul_res1[2087]);
multi_7x28 multi_7x28_mod_2088(clk,rst,matrix_A[2088],matrix_B[88],mul_res1[2088]);
multi_7x28 multi_7x28_mod_2089(clk,rst,matrix_A[2089],matrix_B[89],mul_res1[2089]);
multi_7x28 multi_7x28_mod_2090(clk,rst,matrix_A[2090],matrix_B[90],mul_res1[2090]);
multi_7x28 multi_7x28_mod_2091(clk,rst,matrix_A[2091],matrix_B[91],mul_res1[2091]);
multi_7x28 multi_7x28_mod_2092(clk,rst,matrix_A[2092],matrix_B[92],mul_res1[2092]);
multi_7x28 multi_7x28_mod_2093(clk,rst,matrix_A[2093],matrix_B[93],mul_res1[2093]);
multi_7x28 multi_7x28_mod_2094(clk,rst,matrix_A[2094],matrix_B[94],mul_res1[2094]);
multi_7x28 multi_7x28_mod_2095(clk,rst,matrix_A[2095],matrix_B[95],mul_res1[2095]);
multi_7x28 multi_7x28_mod_2096(clk,rst,matrix_A[2096],matrix_B[96],mul_res1[2096]);
multi_7x28 multi_7x28_mod_2097(clk,rst,matrix_A[2097],matrix_B[97],mul_res1[2097]);
multi_7x28 multi_7x28_mod_2098(clk,rst,matrix_A[2098],matrix_B[98],mul_res1[2098]);
multi_7x28 multi_7x28_mod_2099(clk,rst,matrix_A[2099],matrix_B[99],mul_res1[2099]);
multi_7x28 multi_7x28_mod_2100(clk,rst,matrix_A[2100],matrix_B[100],mul_res1[2100]);
multi_7x28 multi_7x28_mod_2101(clk,rst,matrix_A[2101],matrix_B[101],mul_res1[2101]);
multi_7x28 multi_7x28_mod_2102(clk,rst,matrix_A[2102],matrix_B[102],mul_res1[2102]);
multi_7x28 multi_7x28_mod_2103(clk,rst,matrix_A[2103],matrix_B[103],mul_res1[2103]);
multi_7x28 multi_7x28_mod_2104(clk,rst,matrix_A[2104],matrix_B[104],mul_res1[2104]);
multi_7x28 multi_7x28_mod_2105(clk,rst,matrix_A[2105],matrix_B[105],mul_res1[2105]);
multi_7x28 multi_7x28_mod_2106(clk,rst,matrix_A[2106],matrix_B[106],mul_res1[2106]);
multi_7x28 multi_7x28_mod_2107(clk,rst,matrix_A[2107],matrix_B[107],mul_res1[2107]);
multi_7x28 multi_7x28_mod_2108(clk,rst,matrix_A[2108],matrix_B[108],mul_res1[2108]);
multi_7x28 multi_7x28_mod_2109(clk,rst,matrix_A[2109],matrix_B[109],mul_res1[2109]);
multi_7x28 multi_7x28_mod_2110(clk,rst,matrix_A[2110],matrix_B[110],mul_res1[2110]);
multi_7x28 multi_7x28_mod_2111(clk,rst,matrix_A[2111],matrix_B[111],mul_res1[2111]);
multi_7x28 multi_7x28_mod_2112(clk,rst,matrix_A[2112],matrix_B[112],mul_res1[2112]);
multi_7x28 multi_7x28_mod_2113(clk,rst,matrix_A[2113],matrix_B[113],mul_res1[2113]);
multi_7x28 multi_7x28_mod_2114(clk,rst,matrix_A[2114],matrix_B[114],mul_res1[2114]);
multi_7x28 multi_7x28_mod_2115(clk,rst,matrix_A[2115],matrix_B[115],mul_res1[2115]);
multi_7x28 multi_7x28_mod_2116(clk,rst,matrix_A[2116],matrix_B[116],mul_res1[2116]);
multi_7x28 multi_7x28_mod_2117(clk,rst,matrix_A[2117],matrix_B[117],mul_res1[2117]);
multi_7x28 multi_7x28_mod_2118(clk,rst,matrix_A[2118],matrix_B[118],mul_res1[2118]);
multi_7x28 multi_7x28_mod_2119(clk,rst,matrix_A[2119],matrix_B[119],mul_res1[2119]);
multi_7x28 multi_7x28_mod_2120(clk,rst,matrix_A[2120],matrix_B[120],mul_res1[2120]);
multi_7x28 multi_7x28_mod_2121(clk,rst,matrix_A[2121],matrix_B[121],mul_res1[2121]);
multi_7x28 multi_7x28_mod_2122(clk,rst,matrix_A[2122],matrix_B[122],mul_res1[2122]);
multi_7x28 multi_7x28_mod_2123(clk,rst,matrix_A[2123],matrix_B[123],mul_res1[2123]);
multi_7x28 multi_7x28_mod_2124(clk,rst,matrix_A[2124],matrix_B[124],mul_res1[2124]);
multi_7x28 multi_7x28_mod_2125(clk,rst,matrix_A[2125],matrix_B[125],mul_res1[2125]);
multi_7x28 multi_7x28_mod_2126(clk,rst,matrix_A[2126],matrix_B[126],mul_res1[2126]);
multi_7x28 multi_7x28_mod_2127(clk,rst,matrix_A[2127],matrix_B[127],mul_res1[2127]);
multi_7x28 multi_7x28_mod_2128(clk,rst,matrix_A[2128],matrix_B[128],mul_res1[2128]);
multi_7x28 multi_7x28_mod_2129(clk,rst,matrix_A[2129],matrix_B[129],mul_res1[2129]);
multi_7x28 multi_7x28_mod_2130(clk,rst,matrix_A[2130],matrix_B[130],mul_res1[2130]);
multi_7x28 multi_7x28_mod_2131(clk,rst,matrix_A[2131],matrix_B[131],mul_res1[2131]);
multi_7x28 multi_7x28_mod_2132(clk,rst,matrix_A[2132],matrix_B[132],mul_res1[2132]);
multi_7x28 multi_7x28_mod_2133(clk,rst,matrix_A[2133],matrix_B[133],mul_res1[2133]);
multi_7x28 multi_7x28_mod_2134(clk,rst,matrix_A[2134],matrix_B[134],mul_res1[2134]);
multi_7x28 multi_7x28_mod_2135(clk,rst,matrix_A[2135],matrix_B[135],mul_res1[2135]);
multi_7x28 multi_7x28_mod_2136(clk,rst,matrix_A[2136],matrix_B[136],mul_res1[2136]);
multi_7x28 multi_7x28_mod_2137(clk,rst,matrix_A[2137],matrix_B[137],mul_res1[2137]);
multi_7x28 multi_7x28_mod_2138(clk,rst,matrix_A[2138],matrix_B[138],mul_res1[2138]);
multi_7x28 multi_7x28_mod_2139(clk,rst,matrix_A[2139],matrix_B[139],mul_res1[2139]);
multi_7x28 multi_7x28_mod_2140(clk,rst,matrix_A[2140],matrix_B[140],mul_res1[2140]);
multi_7x28 multi_7x28_mod_2141(clk,rst,matrix_A[2141],matrix_B[141],mul_res1[2141]);
multi_7x28 multi_7x28_mod_2142(clk,rst,matrix_A[2142],matrix_B[142],mul_res1[2142]);
multi_7x28 multi_7x28_mod_2143(clk,rst,matrix_A[2143],matrix_B[143],mul_res1[2143]);
multi_7x28 multi_7x28_mod_2144(clk,rst,matrix_A[2144],matrix_B[144],mul_res1[2144]);
multi_7x28 multi_7x28_mod_2145(clk,rst,matrix_A[2145],matrix_B[145],mul_res1[2145]);
multi_7x28 multi_7x28_mod_2146(clk,rst,matrix_A[2146],matrix_B[146],mul_res1[2146]);
multi_7x28 multi_7x28_mod_2147(clk,rst,matrix_A[2147],matrix_B[147],mul_res1[2147]);
multi_7x28 multi_7x28_mod_2148(clk,rst,matrix_A[2148],matrix_B[148],mul_res1[2148]);
multi_7x28 multi_7x28_mod_2149(clk,rst,matrix_A[2149],matrix_B[149],mul_res1[2149]);
multi_7x28 multi_7x28_mod_2150(clk,rst,matrix_A[2150],matrix_B[150],mul_res1[2150]);
multi_7x28 multi_7x28_mod_2151(clk,rst,matrix_A[2151],matrix_B[151],mul_res1[2151]);
multi_7x28 multi_7x28_mod_2152(clk,rst,matrix_A[2152],matrix_B[152],mul_res1[2152]);
multi_7x28 multi_7x28_mod_2153(clk,rst,matrix_A[2153],matrix_B[153],mul_res1[2153]);
multi_7x28 multi_7x28_mod_2154(clk,rst,matrix_A[2154],matrix_B[154],mul_res1[2154]);
multi_7x28 multi_7x28_mod_2155(clk,rst,matrix_A[2155],matrix_B[155],mul_res1[2155]);
multi_7x28 multi_7x28_mod_2156(clk,rst,matrix_A[2156],matrix_B[156],mul_res1[2156]);
multi_7x28 multi_7x28_mod_2157(clk,rst,matrix_A[2157],matrix_B[157],mul_res1[2157]);
multi_7x28 multi_7x28_mod_2158(clk,rst,matrix_A[2158],matrix_B[158],mul_res1[2158]);
multi_7x28 multi_7x28_mod_2159(clk,rst,matrix_A[2159],matrix_B[159],mul_res1[2159]);
multi_7x28 multi_7x28_mod_2160(clk,rst,matrix_A[2160],matrix_B[160],mul_res1[2160]);
multi_7x28 multi_7x28_mod_2161(clk,rst,matrix_A[2161],matrix_B[161],mul_res1[2161]);
multi_7x28 multi_7x28_mod_2162(clk,rst,matrix_A[2162],matrix_B[162],mul_res1[2162]);
multi_7x28 multi_7x28_mod_2163(clk,rst,matrix_A[2163],matrix_B[163],mul_res1[2163]);
multi_7x28 multi_7x28_mod_2164(clk,rst,matrix_A[2164],matrix_B[164],mul_res1[2164]);
multi_7x28 multi_7x28_mod_2165(clk,rst,matrix_A[2165],matrix_B[165],mul_res1[2165]);
multi_7x28 multi_7x28_mod_2166(clk,rst,matrix_A[2166],matrix_B[166],mul_res1[2166]);
multi_7x28 multi_7x28_mod_2167(clk,rst,matrix_A[2167],matrix_B[167],mul_res1[2167]);
multi_7x28 multi_7x28_mod_2168(clk,rst,matrix_A[2168],matrix_B[168],mul_res1[2168]);
multi_7x28 multi_7x28_mod_2169(clk,rst,matrix_A[2169],matrix_B[169],mul_res1[2169]);
multi_7x28 multi_7x28_mod_2170(clk,rst,matrix_A[2170],matrix_B[170],mul_res1[2170]);
multi_7x28 multi_7x28_mod_2171(clk,rst,matrix_A[2171],matrix_B[171],mul_res1[2171]);
multi_7x28 multi_7x28_mod_2172(clk,rst,matrix_A[2172],matrix_B[172],mul_res1[2172]);
multi_7x28 multi_7x28_mod_2173(clk,rst,matrix_A[2173],matrix_B[173],mul_res1[2173]);
multi_7x28 multi_7x28_mod_2174(clk,rst,matrix_A[2174],matrix_B[174],mul_res1[2174]);
multi_7x28 multi_7x28_mod_2175(clk,rst,matrix_A[2175],matrix_B[175],mul_res1[2175]);
multi_7x28 multi_7x28_mod_2176(clk,rst,matrix_A[2176],matrix_B[176],mul_res1[2176]);
multi_7x28 multi_7x28_mod_2177(clk,rst,matrix_A[2177],matrix_B[177],mul_res1[2177]);
multi_7x28 multi_7x28_mod_2178(clk,rst,matrix_A[2178],matrix_B[178],mul_res1[2178]);
multi_7x28 multi_7x28_mod_2179(clk,rst,matrix_A[2179],matrix_B[179],mul_res1[2179]);
multi_7x28 multi_7x28_mod_2180(clk,rst,matrix_A[2180],matrix_B[180],mul_res1[2180]);
multi_7x28 multi_7x28_mod_2181(clk,rst,matrix_A[2181],matrix_B[181],mul_res1[2181]);
multi_7x28 multi_7x28_mod_2182(clk,rst,matrix_A[2182],matrix_B[182],mul_res1[2182]);
multi_7x28 multi_7x28_mod_2183(clk,rst,matrix_A[2183],matrix_B[183],mul_res1[2183]);
multi_7x28 multi_7x28_mod_2184(clk,rst,matrix_A[2184],matrix_B[184],mul_res1[2184]);
multi_7x28 multi_7x28_mod_2185(clk,rst,matrix_A[2185],matrix_B[185],mul_res1[2185]);
multi_7x28 multi_7x28_mod_2186(clk,rst,matrix_A[2186],matrix_B[186],mul_res1[2186]);
multi_7x28 multi_7x28_mod_2187(clk,rst,matrix_A[2187],matrix_B[187],mul_res1[2187]);
multi_7x28 multi_7x28_mod_2188(clk,rst,matrix_A[2188],matrix_B[188],mul_res1[2188]);
multi_7x28 multi_7x28_mod_2189(clk,rst,matrix_A[2189],matrix_B[189],mul_res1[2189]);
multi_7x28 multi_7x28_mod_2190(clk,rst,matrix_A[2190],matrix_B[190],mul_res1[2190]);
multi_7x28 multi_7x28_mod_2191(clk,rst,matrix_A[2191],matrix_B[191],mul_res1[2191]);
multi_7x28 multi_7x28_mod_2192(clk,rst,matrix_A[2192],matrix_B[192],mul_res1[2192]);
multi_7x28 multi_7x28_mod_2193(clk,rst,matrix_A[2193],matrix_B[193],mul_res1[2193]);
multi_7x28 multi_7x28_mod_2194(clk,rst,matrix_A[2194],matrix_B[194],mul_res1[2194]);
multi_7x28 multi_7x28_mod_2195(clk,rst,matrix_A[2195],matrix_B[195],mul_res1[2195]);
multi_7x28 multi_7x28_mod_2196(clk,rst,matrix_A[2196],matrix_B[196],mul_res1[2196]);
multi_7x28 multi_7x28_mod_2197(clk,rst,matrix_A[2197],matrix_B[197],mul_res1[2197]);
multi_7x28 multi_7x28_mod_2198(clk,rst,matrix_A[2198],matrix_B[198],mul_res1[2198]);
multi_7x28 multi_7x28_mod_2199(clk,rst,matrix_A[2199],matrix_B[199],mul_res1[2199]);
multi_7x28 multi_7x28_mod_2200(clk,rst,matrix_A[2200],matrix_B[0],mul_res1[2200]);
multi_7x28 multi_7x28_mod_2201(clk,rst,matrix_A[2201],matrix_B[1],mul_res1[2201]);
multi_7x28 multi_7x28_mod_2202(clk,rst,matrix_A[2202],matrix_B[2],mul_res1[2202]);
multi_7x28 multi_7x28_mod_2203(clk,rst,matrix_A[2203],matrix_B[3],mul_res1[2203]);
multi_7x28 multi_7x28_mod_2204(clk,rst,matrix_A[2204],matrix_B[4],mul_res1[2204]);
multi_7x28 multi_7x28_mod_2205(clk,rst,matrix_A[2205],matrix_B[5],mul_res1[2205]);
multi_7x28 multi_7x28_mod_2206(clk,rst,matrix_A[2206],matrix_B[6],mul_res1[2206]);
multi_7x28 multi_7x28_mod_2207(clk,rst,matrix_A[2207],matrix_B[7],mul_res1[2207]);
multi_7x28 multi_7x28_mod_2208(clk,rst,matrix_A[2208],matrix_B[8],mul_res1[2208]);
multi_7x28 multi_7x28_mod_2209(clk,rst,matrix_A[2209],matrix_B[9],mul_res1[2209]);
multi_7x28 multi_7x28_mod_2210(clk,rst,matrix_A[2210],matrix_B[10],mul_res1[2210]);
multi_7x28 multi_7x28_mod_2211(clk,rst,matrix_A[2211],matrix_B[11],mul_res1[2211]);
multi_7x28 multi_7x28_mod_2212(clk,rst,matrix_A[2212],matrix_B[12],mul_res1[2212]);
multi_7x28 multi_7x28_mod_2213(clk,rst,matrix_A[2213],matrix_B[13],mul_res1[2213]);
multi_7x28 multi_7x28_mod_2214(clk,rst,matrix_A[2214],matrix_B[14],mul_res1[2214]);
multi_7x28 multi_7x28_mod_2215(clk,rst,matrix_A[2215],matrix_B[15],mul_res1[2215]);
multi_7x28 multi_7x28_mod_2216(clk,rst,matrix_A[2216],matrix_B[16],mul_res1[2216]);
multi_7x28 multi_7x28_mod_2217(clk,rst,matrix_A[2217],matrix_B[17],mul_res1[2217]);
multi_7x28 multi_7x28_mod_2218(clk,rst,matrix_A[2218],matrix_B[18],mul_res1[2218]);
multi_7x28 multi_7x28_mod_2219(clk,rst,matrix_A[2219],matrix_B[19],mul_res1[2219]);
multi_7x28 multi_7x28_mod_2220(clk,rst,matrix_A[2220],matrix_B[20],mul_res1[2220]);
multi_7x28 multi_7x28_mod_2221(clk,rst,matrix_A[2221],matrix_B[21],mul_res1[2221]);
multi_7x28 multi_7x28_mod_2222(clk,rst,matrix_A[2222],matrix_B[22],mul_res1[2222]);
multi_7x28 multi_7x28_mod_2223(clk,rst,matrix_A[2223],matrix_B[23],mul_res1[2223]);
multi_7x28 multi_7x28_mod_2224(clk,rst,matrix_A[2224],matrix_B[24],mul_res1[2224]);
multi_7x28 multi_7x28_mod_2225(clk,rst,matrix_A[2225],matrix_B[25],mul_res1[2225]);
multi_7x28 multi_7x28_mod_2226(clk,rst,matrix_A[2226],matrix_B[26],mul_res1[2226]);
multi_7x28 multi_7x28_mod_2227(clk,rst,matrix_A[2227],matrix_B[27],mul_res1[2227]);
multi_7x28 multi_7x28_mod_2228(clk,rst,matrix_A[2228],matrix_B[28],mul_res1[2228]);
multi_7x28 multi_7x28_mod_2229(clk,rst,matrix_A[2229],matrix_B[29],mul_res1[2229]);
multi_7x28 multi_7x28_mod_2230(clk,rst,matrix_A[2230],matrix_B[30],mul_res1[2230]);
multi_7x28 multi_7x28_mod_2231(clk,rst,matrix_A[2231],matrix_B[31],mul_res1[2231]);
multi_7x28 multi_7x28_mod_2232(clk,rst,matrix_A[2232],matrix_B[32],mul_res1[2232]);
multi_7x28 multi_7x28_mod_2233(clk,rst,matrix_A[2233],matrix_B[33],mul_res1[2233]);
multi_7x28 multi_7x28_mod_2234(clk,rst,matrix_A[2234],matrix_B[34],mul_res1[2234]);
multi_7x28 multi_7x28_mod_2235(clk,rst,matrix_A[2235],matrix_B[35],mul_res1[2235]);
multi_7x28 multi_7x28_mod_2236(clk,rst,matrix_A[2236],matrix_B[36],mul_res1[2236]);
multi_7x28 multi_7x28_mod_2237(clk,rst,matrix_A[2237],matrix_B[37],mul_res1[2237]);
multi_7x28 multi_7x28_mod_2238(clk,rst,matrix_A[2238],matrix_B[38],mul_res1[2238]);
multi_7x28 multi_7x28_mod_2239(clk,rst,matrix_A[2239],matrix_B[39],mul_res1[2239]);
multi_7x28 multi_7x28_mod_2240(clk,rst,matrix_A[2240],matrix_B[40],mul_res1[2240]);
multi_7x28 multi_7x28_mod_2241(clk,rst,matrix_A[2241],matrix_B[41],mul_res1[2241]);
multi_7x28 multi_7x28_mod_2242(clk,rst,matrix_A[2242],matrix_B[42],mul_res1[2242]);
multi_7x28 multi_7x28_mod_2243(clk,rst,matrix_A[2243],matrix_B[43],mul_res1[2243]);
multi_7x28 multi_7x28_mod_2244(clk,rst,matrix_A[2244],matrix_B[44],mul_res1[2244]);
multi_7x28 multi_7x28_mod_2245(clk,rst,matrix_A[2245],matrix_B[45],mul_res1[2245]);
multi_7x28 multi_7x28_mod_2246(clk,rst,matrix_A[2246],matrix_B[46],mul_res1[2246]);
multi_7x28 multi_7x28_mod_2247(clk,rst,matrix_A[2247],matrix_B[47],mul_res1[2247]);
multi_7x28 multi_7x28_mod_2248(clk,rst,matrix_A[2248],matrix_B[48],mul_res1[2248]);
multi_7x28 multi_7x28_mod_2249(clk,rst,matrix_A[2249],matrix_B[49],mul_res1[2249]);
multi_7x28 multi_7x28_mod_2250(clk,rst,matrix_A[2250],matrix_B[50],mul_res1[2250]);
multi_7x28 multi_7x28_mod_2251(clk,rst,matrix_A[2251],matrix_B[51],mul_res1[2251]);
multi_7x28 multi_7x28_mod_2252(clk,rst,matrix_A[2252],matrix_B[52],mul_res1[2252]);
multi_7x28 multi_7x28_mod_2253(clk,rst,matrix_A[2253],matrix_B[53],mul_res1[2253]);
multi_7x28 multi_7x28_mod_2254(clk,rst,matrix_A[2254],matrix_B[54],mul_res1[2254]);
multi_7x28 multi_7x28_mod_2255(clk,rst,matrix_A[2255],matrix_B[55],mul_res1[2255]);
multi_7x28 multi_7x28_mod_2256(clk,rst,matrix_A[2256],matrix_B[56],mul_res1[2256]);
multi_7x28 multi_7x28_mod_2257(clk,rst,matrix_A[2257],matrix_B[57],mul_res1[2257]);
multi_7x28 multi_7x28_mod_2258(clk,rst,matrix_A[2258],matrix_B[58],mul_res1[2258]);
multi_7x28 multi_7x28_mod_2259(clk,rst,matrix_A[2259],matrix_B[59],mul_res1[2259]);
multi_7x28 multi_7x28_mod_2260(clk,rst,matrix_A[2260],matrix_B[60],mul_res1[2260]);
multi_7x28 multi_7x28_mod_2261(clk,rst,matrix_A[2261],matrix_B[61],mul_res1[2261]);
multi_7x28 multi_7x28_mod_2262(clk,rst,matrix_A[2262],matrix_B[62],mul_res1[2262]);
multi_7x28 multi_7x28_mod_2263(clk,rst,matrix_A[2263],matrix_B[63],mul_res1[2263]);
multi_7x28 multi_7x28_mod_2264(clk,rst,matrix_A[2264],matrix_B[64],mul_res1[2264]);
multi_7x28 multi_7x28_mod_2265(clk,rst,matrix_A[2265],matrix_B[65],mul_res1[2265]);
multi_7x28 multi_7x28_mod_2266(clk,rst,matrix_A[2266],matrix_B[66],mul_res1[2266]);
multi_7x28 multi_7x28_mod_2267(clk,rst,matrix_A[2267],matrix_B[67],mul_res1[2267]);
multi_7x28 multi_7x28_mod_2268(clk,rst,matrix_A[2268],matrix_B[68],mul_res1[2268]);
multi_7x28 multi_7x28_mod_2269(clk,rst,matrix_A[2269],matrix_B[69],mul_res1[2269]);
multi_7x28 multi_7x28_mod_2270(clk,rst,matrix_A[2270],matrix_B[70],mul_res1[2270]);
multi_7x28 multi_7x28_mod_2271(clk,rst,matrix_A[2271],matrix_B[71],mul_res1[2271]);
multi_7x28 multi_7x28_mod_2272(clk,rst,matrix_A[2272],matrix_B[72],mul_res1[2272]);
multi_7x28 multi_7x28_mod_2273(clk,rst,matrix_A[2273],matrix_B[73],mul_res1[2273]);
multi_7x28 multi_7x28_mod_2274(clk,rst,matrix_A[2274],matrix_B[74],mul_res1[2274]);
multi_7x28 multi_7x28_mod_2275(clk,rst,matrix_A[2275],matrix_B[75],mul_res1[2275]);
multi_7x28 multi_7x28_mod_2276(clk,rst,matrix_A[2276],matrix_B[76],mul_res1[2276]);
multi_7x28 multi_7x28_mod_2277(clk,rst,matrix_A[2277],matrix_B[77],mul_res1[2277]);
multi_7x28 multi_7x28_mod_2278(clk,rst,matrix_A[2278],matrix_B[78],mul_res1[2278]);
multi_7x28 multi_7x28_mod_2279(clk,rst,matrix_A[2279],matrix_B[79],mul_res1[2279]);
multi_7x28 multi_7x28_mod_2280(clk,rst,matrix_A[2280],matrix_B[80],mul_res1[2280]);
multi_7x28 multi_7x28_mod_2281(clk,rst,matrix_A[2281],matrix_B[81],mul_res1[2281]);
multi_7x28 multi_7x28_mod_2282(clk,rst,matrix_A[2282],matrix_B[82],mul_res1[2282]);
multi_7x28 multi_7x28_mod_2283(clk,rst,matrix_A[2283],matrix_B[83],mul_res1[2283]);
multi_7x28 multi_7x28_mod_2284(clk,rst,matrix_A[2284],matrix_B[84],mul_res1[2284]);
multi_7x28 multi_7x28_mod_2285(clk,rst,matrix_A[2285],matrix_B[85],mul_res1[2285]);
multi_7x28 multi_7x28_mod_2286(clk,rst,matrix_A[2286],matrix_B[86],mul_res1[2286]);
multi_7x28 multi_7x28_mod_2287(clk,rst,matrix_A[2287],matrix_B[87],mul_res1[2287]);
multi_7x28 multi_7x28_mod_2288(clk,rst,matrix_A[2288],matrix_B[88],mul_res1[2288]);
multi_7x28 multi_7x28_mod_2289(clk,rst,matrix_A[2289],matrix_B[89],mul_res1[2289]);
multi_7x28 multi_7x28_mod_2290(clk,rst,matrix_A[2290],matrix_B[90],mul_res1[2290]);
multi_7x28 multi_7x28_mod_2291(clk,rst,matrix_A[2291],matrix_B[91],mul_res1[2291]);
multi_7x28 multi_7x28_mod_2292(clk,rst,matrix_A[2292],matrix_B[92],mul_res1[2292]);
multi_7x28 multi_7x28_mod_2293(clk,rst,matrix_A[2293],matrix_B[93],mul_res1[2293]);
multi_7x28 multi_7x28_mod_2294(clk,rst,matrix_A[2294],matrix_B[94],mul_res1[2294]);
multi_7x28 multi_7x28_mod_2295(clk,rst,matrix_A[2295],matrix_B[95],mul_res1[2295]);
multi_7x28 multi_7x28_mod_2296(clk,rst,matrix_A[2296],matrix_B[96],mul_res1[2296]);
multi_7x28 multi_7x28_mod_2297(clk,rst,matrix_A[2297],matrix_B[97],mul_res1[2297]);
multi_7x28 multi_7x28_mod_2298(clk,rst,matrix_A[2298],matrix_B[98],mul_res1[2298]);
multi_7x28 multi_7x28_mod_2299(clk,rst,matrix_A[2299],matrix_B[99],mul_res1[2299]);
multi_7x28 multi_7x28_mod_2300(clk,rst,matrix_A[2300],matrix_B[100],mul_res1[2300]);
multi_7x28 multi_7x28_mod_2301(clk,rst,matrix_A[2301],matrix_B[101],mul_res1[2301]);
multi_7x28 multi_7x28_mod_2302(clk,rst,matrix_A[2302],matrix_B[102],mul_res1[2302]);
multi_7x28 multi_7x28_mod_2303(clk,rst,matrix_A[2303],matrix_B[103],mul_res1[2303]);
multi_7x28 multi_7x28_mod_2304(clk,rst,matrix_A[2304],matrix_B[104],mul_res1[2304]);
multi_7x28 multi_7x28_mod_2305(clk,rst,matrix_A[2305],matrix_B[105],mul_res1[2305]);
multi_7x28 multi_7x28_mod_2306(clk,rst,matrix_A[2306],matrix_B[106],mul_res1[2306]);
multi_7x28 multi_7x28_mod_2307(clk,rst,matrix_A[2307],matrix_B[107],mul_res1[2307]);
multi_7x28 multi_7x28_mod_2308(clk,rst,matrix_A[2308],matrix_B[108],mul_res1[2308]);
multi_7x28 multi_7x28_mod_2309(clk,rst,matrix_A[2309],matrix_B[109],mul_res1[2309]);
multi_7x28 multi_7x28_mod_2310(clk,rst,matrix_A[2310],matrix_B[110],mul_res1[2310]);
multi_7x28 multi_7x28_mod_2311(clk,rst,matrix_A[2311],matrix_B[111],mul_res1[2311]);
multi_7x28 multi_7x28_mod_2312(clk,rst,matrix_A[2312],matrix_B[112],mul_res1[2312]);
multi_7x28 multi_7x28_mod_2313(clk,rst,matrix_A[2313],matrix_B[113],mul_res1[2313]);
multi_7x28 multi_7x28_mod_2314(clk,rst,matrix_A[2314],matrix_B[114],mul_res1[2314]);
multi_7x28 multi_7x28_mod_2315(clk,rst,matrix_A[2315],matrix_B[115],mul_res1[2315]);
multi_7x28 multi_7x28_mod_2316(clk,rst,matrix_A[2316],matrix_B[116],mul_res1[2316]);
multi_7x28 multi_7x28_mod_2317(clk,rst,matrix_A[2317],matrix_B[117],mul_res1[2317]);
multi_7x28 multi_7x28_mod_2318(clk,rst,matrix_A[2318],matrix_B[118],mul_res1[2318]);
multi_7x28 multi_7x28_mod_2319(clk,rst,matrix_A[2319],matrix_B[119],mul_res1[2319]);
multi_7x28 multi_7x28_mod_2320(clk,rst,matrix_A[2320],matrix_B[120],mul_res1[2320]);
multi_7x28 multi_7x28_mod_2321(clk,rst,matrix_A[2321],matrix_B[121],mul_res1[2321]);
multi_7x28 multi_7x28_mod_2322(clk,rst,matrix_A[2322],matrix_B[122],mul_res1[2322]);
multi_7x28 multi_7x28_mod_2323(clk,rst,matrix_A[2323],matrix_B[123],mul_res1[2323]);
multi_7x28 multi_7x28_mod_2324(clk,rst,matrix_A[2324],matrix_B[124],mul_res1[2324]);
multi_7x28 multi_7x28_mod_2325(clk,rst,matrix_A[2325],matrix_B[125],mul_res1[2325]);
multi_7x28 multi_7x28_mod_2326(clk,rst,matrix_A[2326],matrix_B[126],mul_res1[2326]);
multi_7x28 multi_7x28_mod_2327(clk,rst,matrix_A[2327],matrix_B[127],mul_res1[2327]);
multi_7x28 multi_7x28_mod_2328(clk,rst,matrix_A[2328],matrix_B[128],mul_res1[2328]);
multi_7x28 multi_7x28_mod_2329(clk,rst,matrix_A[2329],matrix_B[129],mul_res1[2329]);
multi_7x28 multi_7x28_mod_2330(clk,rst,matrix_A[2330],matrix_B[130],mul_res1[2330]);
multi_7x28 multi_7x28_mod_2331(clk,rst,matrix_A[2331],matrix_B[131],mul_res1[2331]);
multi_7x28 multi_7x28_mod_2332(clk,rst,matrix_A[2332],matrix_B[132],mul_res1[2332]);
multi_7x28 multi_7x28_mod_2333(clk,rst,matrix_A[2333],matrix_B[133],mul_res1[2333]);
multi_7x28 multi_7x28_mod_2334(clk,rst,matrix_A[2334],matrix_B[134],mul_res1[2334]);
multi_7x28 multi_7x28_mod_2335(clk,rst,matrix_A[2335],matrix_B[135],mul_res1[2335]);
multi_7x28 multi_7x28_mod_2336(clk,rst,matrix_A[2336],matrix_B[136],mul_res1[2336]);
multi_7x28 multi_7x28_mod_2337(clk,rst,matrix_A[2337],matrix_B[137],mul_res1[2337]);
multi_7x28 multi_7x28_mod_2338(clk,rst,matrix_A[2338],matrix_B[138],mul_res1[2338]);
multi_7x28 multi_7x28_mod_2339(clk,rst,matrix_A[2339],matrix_B[139],mul_res1[2339]);
multi_7x28 multi_7x28_mod_2340(clk,rst,matrix_A[2340],matrix_B[140],mul_res1[2340]);
multi_7x28 multi_7x28_mod_2341(clk,rst,matrix_A[2341],matrix_B[141],mul_res1[2341]);
multi_7x28 multi_7x28_mod_2342(clk,rst,matrix_A[2342],matrix_B[142],mul_res1[2342]);
multi_7x28 multi_7x28_mod_2343(clk,rst,matrix_A[2343],matrix_B[143],mul_res1[2343]);
multi_7x28 multi_7x28_mod_2344(clk,rst,matrix_A[2344],matrix_B[144],mul_res1[2344]);
multi_7x28 multi_7x28_mod_2345(clk,rst,matrix_A[2345],matrix_B[145],mul_res1[2345]);
multi_7x28 multi_7x28_mod_2346(clk,rst,matrix_A[2346],matrix_B[146],mul_res1[2346]);
multi_7x28 multi_7x28_mod_2347(clk,rst,matrix_A[2347],matrix_B[147],mul_res1[2347]);
multi_7x28 multi_7x28_mod_2348(clk,rst,matrix_A[2348],matrix_B[148],mul_res1[2348]);
multi_7x28 multi_7x28_mod_2349(clk,rst,matrix_A[2349],matrix_B[149],mul_res1[2349]);
multi_7x28 multi_7x28_mod_2350(clk,rst,matrix_A[2350],matrix_B[150],mul_res1[2350]);
multi_7x28 multi_7x28_mod_2351(clk,rst,matrix_A[2351],matrix_B[151],mul_res1[2351]);
multi_7x28 multi_7x28_mod_2352(clk,rst,matrix_A[2352],matrix_B[152],mul_res1[2352]);
multi_7x28 multi_7x28_mod_2353(clk,rst,matrix_A[2353],matrix_B[153],mul_res1[2353]);
multi_7x28 multi_7x28_mod_2354(clk,rst,matrix_A[2354],matrix_B[154],mul_res1[2354]);
multi_7x28 multi_7x28_mod_2355(clk,rst,matrix_A[2355],matrix_B[155],mul_res1[2355]);
multi_7x28 multi_7x28_mod_2356(clk,rst,matrix_A[2356],matrix_B[156],mul_res1[2356]);
multi_7x28 multi_7x28_mod_2357(clk,rst,matrix_A[2357],matrix_B[157],mul_res1[2357]);
multi_7x28 multi_7x28_mod_2358(clk,rst,matrix_A[2358],matrix_B[158],mul_res1[2358]);
multi_7x28 multi_7x28_mod_2359(clk,rst,matrix_A[2359],matrix_B[159],mul_res1[2359]);
multi_7x28 multi_7x28_mod_2360(clk,rst,matrix_A[2360],matrix_B[160],mul_res1[2360]);
multi_7x28 multi_7x28_mod_2361(clk,rst,matrix_A[2361],matrix_B[161],mul_res1[2361]);
multi_7x28 multi_7x28_mod_2362(clk,rst,matrix_A[2362],matrix_B[162],mul_res1[2362]);
multi_7x28 multi_7x28_mod_2363(clk,rst,matrix_A[2363],matrix_B[163],mul_res1[2363]);
multi_7x28 multi_7x28_mod_2364(clk,rst,matrix_A[2364],matrix_B[164],mul_res1[2364]);
multi_7x28 multi_7x28_mod_2365(clk,rst,matrix_A[2365],matrix_B[165],mul_res1[2365]);
multi_7x28 multi_7x28_mod_2366(clk,rst,matrix_A[2366],matrix_B[166],mul_res1[2366]);
multi_7x28 multi_7x28_mod_2367(clk,rst,matrix_A[2367],matrix_B[167],mul_res1[2367]);
multi_7x28 multi_7x28_mod_2368(clk,rst,matrix_A[2368],matrix_B[168],mul_res1[2368]);
multi_7x28 multi_7x28_mod_2369(clk,rst,matrix_A[2369],matrix_B[169],mul_res1[2369]);
multi_7x28 multi_7x28_mod_2370(clk,rst,matrix_A[2370],matrix_B[170],mul_res1[2370]);
multi_7x28 multi_7x28_mod_2371(clk,rst,matrix_A[2371],matrix_B[171],mul_res1[2371]);
multi_7x28 multi_7x28_mod_2372(clk,rst,matrix_A[2372],matrix_B[172],mul_res1[2372]);
multi_7x28 multi_7x28_mod_2373(clk,rst,matrix_A[2373],matrix_B[173],mul_res1[2373]);
multi_7x28 multi_7x28_mod_2374(clk,rst,matrix_A[2374],matrix_B[174],mul_res1[2374]);
multi_7x28 multi_7x28_mod_2375(clk,rst,matrix_A[2375],matrix_B[175],mul_res1[2375]);
multi_7x28 multi_7x28_mod_2376(clk,rst,matrix_A[2376],matrix_B[176],mul_res1[2376]);
multi_7x28 multi_7x28_mod_2377(clk,rst,matrix_A[2377],matrix_B[177],mul_res1[2377]);
multi_7x28 multi_7x28_mod_2378(clk,rst,matrix_A[2378],matrix_B[178],mul_res1[2378]);
multi_7x28 multi_7x28_mod_2379(clk,rst,matrix_A[2379],matrix_B[179],mul_res1[2379]);
multi_7x28 multi_7x28_mod_2380(clk,rst,matrix_A[2380],matrix_B[180],mul_res1[2380]);
multi_7x28 multi_7x28_mod_2381(clk,rst,matrix_A[2381],matrix_B[181],mul_res1[2381]);
multi_7x28 multi_7x28_mod_2382(clk,rst,matrix_A[2382],matrix_B[182],mul_res1[2382]);
multi_7x28 multi_7x28_mod_2383(clk,rst,matrix_A[2383],matrix_B[183],mul_res1[2383]);
multi_7x28 multi_7x28_mod_2384(clk,rst,matrix_A[2384],matrix_B[184],mul_res1[2384]);
multi_7x28 multi_7x28_mod_2385(clk,rst,matrix_A[2385],matrix_B[185],mul_res1[2385]);
multi_7x28 multi_7x28_mod_2386(clk,rst,matrix_A[2386],matrix_B[186],mul_res1[2386]);
multi_7x28 multi_7x28_mod_2387(clk,rst,matrix_A[2387],matrix_B[187],mul_res1[2387]);
multi_7x28 multi_7x28_mod_2388(clk,rst,matrix_A[2388],matrix_B[188],mul_res1[2388]);
multi_7x28 multi_7x28_mod_2389(clk,rst,matrix_A[2389],matrix_B[189],mul_res1[2389]);
multi_7x28 multi_7x28_mod_2390(clk,rst,matrix_A[2390],matrix_B[190],mul_res1[2390]);
multi_7x28 multi_7x28_mod_2391(clk,rst,matrix_A[2391],matrix_B[191],mul_res1[2391]);
multi_7x28 multi_7x28_mod_2392(clk,rst,matrix_A[2392],matrix_B[192],mul_res1[2392]);
multi_7x28 multi_7x28_mod_2393(clk,rst,matrix_A[2393],matrix_B[193],mul_res1[2393]);
multi_7x28 multi_7x28_mod_2394(clk,rst,matrix_A[2394],matrix_B[194],mul_res1[2394]);
multi_7x28 multi_7x28_mod_2395(clk,rst,matrix_A[2395],matrix_B[195],mul_res1[2395]);
multi_7x28 multi_7x28_mod_2396(clk,rst,matrix_A[2396],matrix_B[196],mul_res1[2396]);
multi_7x28 multi_7x28_mod_2397(clk,rst,matrix_A[2397],matrix_B[197],mul_res1[2397]);
multi_7x28 multi_7x28_mod_2398(clk,rst,matrix_A[2398],matrix_B[198],mul_res1[2398]);
multi_7x28 multi_7x28_mod_2399(clk,rst,matrix_A[2399],matrix_B[199],mul_res1[2399]);
multi_7x28 multi_7x28_mod_2400(clk,rst,matrix_A[2400],matrix_B[0],mul_res1[2400]);
multi_7x28 multi_7x28_mod_2401(clk,rst,matrix_A[2401],matrix_B[1],mul_res1[2401]);
multi_7x28 multi_7x28_mod_2402(clk,rst,matrix_A[2402],matrix_B[2],mul_res1[2402]);
multi_7x28 multi_7x28_mod_2403(clk,rst,matrix_A[2403],matrix_B[3],mul_res1[2403]);
multi_7x28 multi_7x28_mod_2404(clk,rst,matrix_A[2404],matrix_B[4],mul_res1[2404]);
multi_7x28 multi_7x28_mod_2405(clk,rst,matrix_A[2405],matrix_B[5],mul_res1[2405]);
multi_7x28 multi_7x28_mod_2406(clk,rst,matrix_A[2406],matrix_B[6],mul_res1[2406]);
multi_7x28 multi_7x28_mod_2407(clk,rst,matrix_A[2407],matrix_B[7],mul_res1[2407]);
multi_7x28 multi_7x28_mod_2408(clk,rst,matrix_A[2408],matrix_B[8],mul_res1[2408]);
multi_7x28 multi_7x28_mod_2409(clk,rst,matrix_A[2409],matrix_B[9],mul_res1[2409]);
multi_7x28 multi_7x28_mod_2410(clk,rst,matrix_A[2410],matrix_B[10],mul_res1[2410]);
multi_7x28 multi_7x28_mod_2411(clk,rst,matrix_A[2411],matrix_B[11],mul_res1[2411]);
multi_7x28 multi_7x28_mod_2412(clk,rst,matrix_A[2412],matrix_B[12],mul_res1[2412]);
multi_7x28 multi_7x28_mod_2413(clk,rst,matrix_A[2413],matrix_B[13],mul_res1[2413]);
multi_7x28 multi_7x28_mod_2414(clk,rst,matrix_A[2414],matrix_B[14],mul_res1[2414]);
multi_7x28 multi_7x28_mod_2415(clk,rst,matrix_A[2415],matrix_B[15],mul_res1[2415]);
multi_7x28 multi_7x28_mod_2416(clk,rst,matrix_A[2416],matrix_B[16],mul_res1[2416]);
multi_7x28 multi_7x28_mod_2417(clk,rst,matrix_A[2417],matrix_B[17],mul_res1[2417]);
multi_7x28 multi_7x28_mod_2418(clk,rst,matrix_A[2418],matrix_B[18],mul_res1[2418]);
multi_7x28 multi_7x28_mod_2419(clk,rst,matrix_A[2419],matrix_B[19],mul_res1[2419]);
multi_7x28 multi_7x28_mod_2420(clk,rst,matrix_A[2420],matrix_B[20],mul_res1[2420]);
multi_7x28 multi_7x28_mod_2421(clk,rst,matrix_A[2421],matrix_B[21],mul_res1[2421]);
multi_7x28 multi_7x28_mod_2422(clk,rst,matrix_A[2422],matrix_B[22],mul_res1[2422]);
multi_7x28 multi_7x28_mod_2423(clk,rst,matrix_A[2423],matrix_B[23],mul_res1[2423]);
multi_7x28 multi_7x28_mod_2424(clk,rst,matrix_A[2424],matrix_B[24],mul_res1[2424]);
multi_7x28 multi_7x28_mod_2425(clk,rst,matrix_A[2425],matrix_B[25],mul_res1[2425]);
multi_7x28 multi_7x28_mod_2426(clk,rst,matrix_A[2426],matrix_B[26],mul_res1[2426]);
multi_7x28 multi_7x28_mod_2427(clk,rst,matrix_A[2427],matrix_B[27],mul_res1[2427]);
multi_7x28 multi_7x28_mod_2428(clk,rst,matrix_A[2428],matrix_B[28],mul_res1[2428]);
multi_7x28 multi_7x28_mod_2429(clk,rst,matrix_A[2429],matrix_B[29],mul_res1[2429]);
multi_7x28 multi_7x28_mod_2430(clk,rst,matrix_A[2430],matrix_B[30],mul_res1[2430]);
multi_7x28 multi_7x28_mod_2431(clk,rst,matrix_A[2431],matrix_B[31],mul_res1[2431]);
multi_7x28 multi_7x28_mod_2432(clk,rst,matrix_A[2432],matrix_B[32],mul_res1[2432]);
multi_7x28 multi_7x28_mod_2433(clk,rst,matrix_A[2433],matrix_B[33],mul_res1[2433]);
multi_7x28 multi_7x28_mod_2434(clk,rst,matrix_A[2434],matrix_B[34],mul_res1[2434]);
multi_7x28 multi_7x28_mod_2435(clk,rst,matrix_A[2435],matrix_B[35],mul_res1[2435]);
multi_7x28 multi_7x28_mod_2436(clk,rst,matrix_A[2436],matrix_B[36],mul_res1[2436]);
multi_7x28 multi_7x28_mod_2437(clk,rst,matrix_A[2437],matrix_B[37],mul_res1[2437]);
multi_7x28 multi_7x28_mod_2438(clk,rst,matrix_A[2438],matrix_B[38],mul_res1[2438]);
multi_7x28 multi_7x28_mod_2439(clk,rst,matrix_A[2439],matrix_B[39],mul_res1[2439]);
multi_7x28 multi_7x28_mod_2440(clk,rst,matrix_A[2440],matrix_B[40],mul_res1[2440]);
multi_7x28 multi_7x28_mod_2441(clk,rst,matrix_A[2441],matrix_B[41],mul_res1[2441]);
multi_7x28 multi_7x28_mod_2442(clk,rst,matrix_A[2442],matrix_B[42],mul_res1[2442]);
multi_7x28 multi_7x28_mod_2443(clk,rst,matrix_A[2443],matrix_B[43],mul_res1[2443]);
multi_7x28 multi_7x28_mod_2444(clk,rst,matrix_A[2444],matrix_B[44],mul_res1[2444]);
multi_7x28 multi_7x28_mod_2445(clk,rst,matrix_A[2445],matrix_B[45],mul_res1[2445]);
multi_7x28 multi_7x28_mod_2446(clk,rst,matrix_A[2446],matrix_B[46],mul_res1[2446]);
multi_7x28 multi_7x28_mod_2447(clk,rst,matrix_A[2447],matrix_B[47],mul_res1[2447]);
multi_7x28 multi_7x28_mod_2448(clk,rst,matrix_A[2448],matrix_B[48],mul_res1[2448]);
multi_7x28 multi_7x28_mod_2449(clk,rst,matrix_A[2449],matrix_B[49],mul_res1[2449]);
multi_7x28 multi_7x28_mod_2450(clk,rst,matrix_A[2450],matrix_B[50],mul_res1[2450]);
multi_7x28 multi_7x28_mod_2451(clk,rst,matrix_A[2451],matrix_B[51],mul_res1[2451]);
multi_7x28 multi_7x28_mod_2452(clk,rst,matrix_A[2452],matrix_B[52],mul_res1[2452]);
multi_7x28 multi_7x28_mod_2453(clk,rst,matrix_A[2453],matrix_B[53],mul_res1[2453]);
multi_7x28 multi_7x28_mod_2454(clk,rst,matrix_A[2454],matrix_B[54],mul_res1[2454]);
multi_7x28 multi_7x28_mod_2455(clk,rst,matrix_A[2455],matrix_B[55],mul_res1[2455]);
multi_7x28 multi_7x28_mod_2456(clk,rst,matrix_A[2456],matrix_B[56],mul_res1[2456]);
multi_7x28 multi_7x28_mod_2457(clk,rst,matrix_A[2457],matrix_B[57],mul_res1[2457]);
multi_7x28 multi_7x28_mod_2458(clk,rst,matrix_A[2458],matrix_B[58],mul_res1[2458]);
multi_7x28 multi_7x28_mod_2459(clk,rst,matrix_A[2459],matrix_B[59],mul_res1[2459]);
multi_7x28 multi_7x28_mod_2460(clk,rst,matrix_A[2460],matrix_B[60],mul_res1[2460]);
multi_7x28 multi_7x28_mod_2461(clk,rst,matrix_A[2461],matrix_B[61],mul_res1[2461]);
multi_7x28 multi_7x28_mod_2462(clk,rst,matrix_A[2462],matrix_B[62],mul_res1[2462]);
multi_7x28 multi_7x28_mod_2463(clk,rst,matrix_A[2463],matrix_B[63],mul_res1[2463]);
multi_7x28 multi_7x28_mod_2464(clk,rst,matrix_A[2464],matrix_B[64],mul_res1[2464]);
multi_7x28 multi_7x28_mod_2465(clk,rst,matrix_A[2465],matrix_B[65],mul_res1[2465]);
multi_7x28 multi_7x28_mod_2466(clk,rst,matrix_A[2466],matrix_B[66],mul_res1[2466]);
multi_7x28 multi_7x28_mod_2467(clk,rst,matrix_A[2467],matrix_B[67],mul_res1[2467]);
multi_7x28 multi_7x28_mod_2468(clk,rst,matrix_A[2468],matrix_B[68],mul_res1[2468]);
multi_7x28 multi_7x28_mod_2469(clk,rst,matrix_A[2469],matrix_B[69],mul_res1[2469]);
multi_7x28 multi_7x28_mod_2470(clk,rst,matrix_A[2470],matrix_B[70],mul_res1[2470]);
multi_7x28 multi_7x28_mod_2471(clk,rst,matrix_A[2471],matrix_B[71],mul_res1[2471]);
multi_7x28 multi_7x28_mod_2472(clk,rst,matrix_A[2472],matrix_B[72],mul_res1[2472]);
multi_7x28 multi_7x28_mod_2473(clk,rst,matrix_A[2473],matrix_B[73],mul_res1[2473]);
multi_7x28 multi_7x28_mod_2474(clk,rst,matrix_A[2474],matrix_B[74],mul_res1[2474]);
multi_7x28 multi_7x28_mod_2475(clk,rst,matrix_A[2475],matrix_B[75],mul_res1[2475]);
multi_7x28 multi_7x28_mod_2476(clk,rst,matrix_A[2476],matrix_B[76],mul_res1[2476]);
multi_7x28 multi_7x28_mod_2477(clk,rst,matrix_A[2477],matrix_B[77],mul_res1[2477]);
multi_7x28 multi_7x28_mod_2478(clk,rst,matrix_A[2478],matrix_B[78],mul_res1[2478]);
multi_7x28 multi_7x28_mod_2479(clk,rst,matrix_A[2479],matrix_B[79],mul_res1[2479]);
multi_7x28 multi_7x28_mod_2480(clk,rst,matrix_A[2480],matrix_B[80],mul_res1[2480]);
multi_7x28 multi_7x28_mod_2481(clk,rst,matrix_A[2481],matrix_B[81],mul_res1[2481]);
multi_7x28 multi_7x28_mod_2482(clk,rst,matrix_A[2482],matrix_B[82],mul_res1[2482]);
multi_7x28 multi_7x28_mod_2483(clk,rst,matrix_A[2483],matrix_B[83],mul_res1[2483]);
multi_7x28 multi_7x28_mod_2484(clk,rst,matrix_A[2484],matrix_B[84],mul_res1[2484]);
multi_7x28 multi_7x28_mod_2485(clk,rst,matrix_A[2485],matrix_B[85],mul_res1[2485]);
multi_7x28 multi_7x28_mod_2486(clk,rst,matrix_A[2486],matrix_B[86],mul_res1[2486]);
multi_7x28 multi_7x28_mod_2487(clk,rst,matrix_A[2487],matrix_B[87],mul_res1[2487]);
multi_7x28 multi_7x28_mod_2488(clk,rst,matrix_A[2488],matrix_B[88],mul_res1[2488]);
multi_7x28 multi_7x28_mod_2489(clk,rst,matrix_A[2489],matrix_B[89],mul_res1[2489]);
multi_7x28 multi_7x28_mod_2490(clk,rst,matrix_A[2490],matrix_B[90],mul_res1[2490]);
multi_7x28 multi_7x28_mod_2491(clk,rst,matrix_A[2491],matrix_B[91],mul_res1[2491]);
multi_7x28 multi_7x28_mod_2492(clk,rst,matrix_A[2492],matrix_B[92],mul_res1[2492]);
multi_7x28 multi_7x28_mod_2493(clk,rst,matrix_A[2493],matrix_B[93],mul_res1[2493]);
multi_7x28 multi_7x28_mod_2494(clk,rst,matrix_A[2494],matrix_B[94],mul_res1[2494]);
multi_7x28 multi_7x28_mod_2495(clk,rst,matrix_A[2495],matrix_B[95],mul_res1[2495]);
multi_7x28 multi_7x28_mod_2496(clk,rst,matrix_A[2496],matrix_B[96],mul_res1[2496]);
multi_7x28 multi_7x28_mod_2497(clk,rst,matrix_A[2497],matrix_B[97],mul_res1[2497]);
multi_7x28 multi_7x28_mod_2498(clk,rst,matrix_A[2498],matrix_B[98],mul_res1[2498]);
multi_7x28 multi_7x28_mod_2499(clk,rst,matrix_A[2499],matrix_B[99],mul_res1[2499]);
multi_7x28 multi_7x28_mod_2500(clk,rst,matrix_A[2500],matrix_B[100],mul_res1[2500]);
multi_7x28 multi_7x28_mod_2501(clk,rst,matrix_A[2501],matrix_B[101],mul_res1[2501]);
multi_7x28 multi_7x28_mod_2502(clk,rst,matrix_A[2502],matrix_B[102],mul_res1[2502]);
multi_7x28 multi_7x28_mod_2503(clk,rst,matrix_A[2503],matrix_B[103],mul_res1[2503]);
multi_7x28 multi_7x28_mod_2504(clk,rst,matrix_A[2504],matrix_B[104],mul_res1[2504]);
multi_7x28 multi_7x28_mod_2505(clk,rst,matrix_A[2505],matrix_B[105],mul_res1[2505]);
multi_7x28 multi_7x28_mod_2506(clk,rst,matrix_A[2506],matrix_B[106],mul_res1[2506]);
multi_7x28 multi_7x28_mod_2507(clk,rst,matrix_A[2507],matrix_B[107],mul_res1[2507]);
multi_7x28 multi_7x28_mod_2508(clk,rst,matrix_A[2508],matrix_B[108],mul_res1[2508]);
multi_7x28 multi_7x28_mod_2509(clk,rst,matrix_A[2509],matrix_B[109],mul_res1[2509]);
multi_7x28 multi_7x28_mod_2510(clk,rst,matrix_A[2510],matrix_B[110],mul_res1[2510]);
multi_7x28 multi_7x28_mod_2511(clk,rst,matrix_A[2511],matrix_B[111],mul_res1[2511]);
multi_7x28 multi_7x28_mod_2512(clk,rst,matrix_A[2512],matrix_B[112],mul_res1[2512]);
multi_7x28 multi_7x28_mod_2513(clk,rst,matrix_A[2513],matrix_B[113],mul_res1[2513]);
multi_7x28 multi_7x28_mod_2514(clk,rst,matrix_A[2514],matrix_B[114],mul_res1[2514]);
multi_7x28 multi_7x28_mod_2515(clk,rst,matrix_A[2515],matrix_B[115],mul_res1[2515]);
multi_7x28 multi_7x28_mod_2516(clk,rst,matrix_A[2516],matrix_B[116],mul_res1[2516]);
multi_7x28 multi_7x28_mod_2517(clk,rst,matrix_A[2517],matrix_B[117],mul_res1[2517]);
multi_7x28 multi_7x28_mod_2518(clk,rst,matrix_A[2518],matrix_B[118],mul_res1[2518]);
multi_7x28 multi_7x28_mod_2519(clk,rst,matrix_A[2519],matrix_B[119],mul_res1[2519]);
multi_7x28 multi_7x28_mod_2520(clk,rst,matrix_A[2520],matrix_B[120],mul_res1[2520]);
multi_7x28 multi_7x28_mod_2521(clk,rst,matrix_A[2521],matrix_B[121],mul_res1[2521]);
multi_7x28 multi_7x28_mod_2522(clk,rst,matrix_A[2522],matrix_B[122],mul_res1[2522]);
multi_7x28 multi_7x28_mod_2523(clk,rst,matrix_A[2523],matrix_B[123],mul_res1[2523]);
multi_7x28 multi_7x28_mod_2524(clk,rst,matrix_A[2524],matrix_B[124],mul_res1[2524]);
multi_7x28 multi_7x28_mod_2525(clk,rst,matrix_A[2525],matrix_B[125],mul_res1[2525]);
multi_7x28 multi_7x28_mod_2526(clk,rst,matrix_A[2526],matrix_B[126],mul_res1[2526]);
multi_7x28 multi_7x28_mod_2527(clk,rst,matrix_A[2527],matrix_B[127],mul_res1[2527]);
multi_7x28 multi_7x28_mod_2528(clk,rst,matrix_A[2528],matrix_B[128],mul_res1[2528]);
multi_7x28 multi_7x28_mod_2529(clk,rst,matrix_A[2529],matrix_B[129],mul_res1[2529]);
multi_7x28 multi_7x28_mod_2530(clk,rst,matrix_A[2530],matrix_B[130],mul_res1[2530]);
multi_7x28 multi_7x28_mod_2531(clk,rst,matrix_A[2531],matrix_B[131],mul_res1[2531]);
multi_7x28 multi_7x28_mod_2532(clk,rst,matrix_A[2532],matrix_B[132],mul_res1[2532]);
multi_7x28 multi_7x28_mod_2533(clk,rst,matrix_A[2533],matrix_B[133],mul_res1[2533]);
multi_7x28 multi_7x28_mod_2534(clk,rst,matrix_A[2534],matrix_B[134],mul_res1[2534]);
multi_7x28 multi_7x28_mod_2535(clk,rst,matrix_A[2535],matrix_B[135],mul_res1[2535]);
multi_7x28 multi_7x28_mod_2536(clk,rst,matrix_A[2536],matrix_B[136],mul_res1[2536]);
multi_7x28 multi_7x28_mod_2537(clk,rst,matrix_A[2537],matrix_B[137],mul_res1[2537]);
multi_7x28 multi_7x28_mod_2538(clk,rst,matrix_A[2538],matrix_B[138],mul_res1[2538]);
multi_7x28 multi_7x28_mod_2539(clk,rst,matrix_A[2539],matrix_B[139],mul_res1[2539]);
multi_7x28 multi_7x28_mod_2540(clk,rst,matrix_A[2540],matrix_B[140],mul_res1[2540]);
multi_7x28 multi_7x28_mod_2541(clk,rst,matrix_A[2541],matrix_B[141],mul_res1[2541]);
multi_7x28 multi_7x28_mod_2542(clk,rst,matrix_A[2542],matrix_B[142],mul_res1[2542]);
multi_7x28 multi_7x28_mod_2543(clk,rst,matrix_A[2543],matrix_B[143],mul_res1[2543]);
multi_7x28 multi_7x28_mod_2544(clk,rst,matrix_A[2544],matrix_B[144],mul_res1[2544]);
multi_7x28 multi_7x28_mod_2545(clk,rst,matrix_A[2545],matrix_B[145],mul_res1[2545]);
multi_7x28 multi_7x28_mod_2546(clk,rst,matrix_A[2546],matrix_B[146],mul_res1[2546]);
multi_7x28 multi_7x28_mod_2547(clk,rst,matrix_A[2547],matrix_B[147],mul_res1[2547]);
multi_7x28 multi_7x28_mod_2548(clk,rst,matrix_A[2548],matrix_B[148],mul_res1[2548]);
multi_7x28 multi_7x28_mod_2549(clk,rst,matrix_A[2549],matrix_B[149],mul_res1[2549]);
multi_7x28 multi_7x28_mod_2550(clk,rst,matrix_A[2550],matrix_B[150],mul_res1[2550]);
multi_7x28 multi_7x28_mod_2551(clk,rst,matrix_A[2551],matrix_B[151],mul_res1[2551]);
multi_7x28 multi_7x28_mod_2552(clk,rst,matrix_A[2552],matrix_B[152],mul_res1[2552]);
multi_7x28 multi_7x28_mod_2553(clk,rst,matrix_A[2553],matrix_B[153],mul_res1[2553]);
multi_7x28 multi_7x28_mod_2554(clk,rst,matrix_A[2554],matrix_B[154],mul_res1[2554]);
multi_7x28 multi_7x28_mod_2555(clk,rst,matrix_A[2555],matrix_B[155],mul_res1[2555]);
multi_7x28 multi_7x28_mod_2556(clk,rst,matrix_A[2556],matrix_B[156],mul_res1[2556]);
multi_7x28 multi_7x28_mod_2557(clk,rst,matrix_A[2557],matrix_B[157],mul_res1[2557]);
multi_7x28 multi_7x28_mod_2558(clk,rst,matrix_A[2558],matrix_B[158],mul_res1[2558]);
multi_7x28 multi_7x28_mod_2559(clk,rst,matrix_A[2559],matrix_B[159],mul_res1[2559]);
multi_7x28 multi_7x28_mod_2560(clk,rst,matrix_A[2560],matrix_B[160],mul_res1[2560]);
multi_7x28 multi_7x28_mod_2561(clk,rst,matrix_A[2561],matrix_B[161],mul_res1[2561]);
multi_7x28 multi_7x28_mod_2562(clk,rst,matrix_A[2562],matrix_B[162],mul_res1[2562]);
multi_7x28 multi_7x28_mod_2563(clk,rst,matrix_A[2563],matrix_B[163],mul_res1[2563]);
multi_7x28 multi_7x28_mod_2564(clk,rst,matrix_A[2564],matrix_B[164],mul_res1[2564]);
multi_7x28 multi_7x28_mod_2565(clk,rst,matrix_A[2565],matrix_B[165],mul_res1[2565]);
multi_7x28 multi_7x28_mod_2566(clk,rst,matrix_A[2566],matrix_B[166],mul_res1[2566]);
multi_7x28 multi_7x28_mod_2567(clk,rst,matrix_A[2567],matrix_B[167],mul_res1[2567]);
multi_7x28 multi_7x28_mod_2568(clk,rst,matrix_A[2568],matrix_B[168],mul_res1[2568]);
multi_7x28 multi_7x28_mod_2569(clk,rst,matrix_A[2569],matrix_B[169],mul_res1[2569]);
multi_7x28 multi_7x28_mod_2570(clk,rst,matrix_A[2570],matrix_B[170],mul_res1[2570]);
multi_7x28 multi_7x28_mod_2571(clk,rst,matrix_A[2571],matrix_B[171],mul_res1[2571]);
multi_7x28 multi_7x28_mod_2572(clk,rst,matrix_A[2572],matrix_B[172],mul_res1[2572]);
multi_7x28 multi_7x28_mod_2573(clk,rst,matrix_A[2573],matrix_B[173],mul_res1[2573]);
multi_7x28 multi_7x28_mod_2574(clk,rst,matrix_A[2574],matrix_B[174],mul_res1[2574]);
multi_7x28 multi_7x28_mod_2575(clk,rst,matrix_A[2575],matrix_B[175],mul_res1[2575]);
multi_7x28 multi_7x28_mod_2576(clk,rst,matrix_A[2576],matrix_B[176],mul_res1[2576]);
multi_7x28 multi_7x28_mod_2577(clk,rst,matrix_A[2577],matrix_B[177],mul_res1[2577]);
multi_7x28 multi_7x28_mod_2578(clk,rst,matrix_A[2578],matrix_B[178],mul_res1[2578]);
multi_7x28 multi_7x28_mod_2579(clk,rst,matrix_A[2579],matrix_B[179],mul_res1[2579]);
multi_7x28 multi_7x28_mod_2580(clk,rst,matrix_A[2580],matrix_B[180],mul_res1[2580]);
multi_7x28 multi_7x28_mod_2581(clk,rst,matrix_A[2581],matrix_B[181],mul_res1[2581]);
multi_7x28 multi_7x28_mod_2582(clk,rst,matrix_A[2582],matrix_B[182],mul_res1[2582]);
multi_7x28 multi_7x28_mod_2583(clk,rst,matrix_A[2583],matrix_B[183],mul_res1[2583]);
multi_7x28 multi_7x28_mod_2584(clk,rst,matrix_A[2584],matrix_B[184],mul_res1[2584]);
multi_7x28 multi_7x28_mod_2585(clk,rst,matrix_A[2585],matrix_B[185],mul_res1[2585]);
multi_7x28 multi_7x28_mod_2586(clk,rst,matrix_A[2586],matrix_B[186],mul_res1[2586]);
multi_7x28 multi_7x28_mod_2587(clk,rst,matrix_A[2587],matrix_B[187],mul_res1[2587]);
multi_7x28 multi_7x28_mod_2588(clk,rst,matrix_A[2588],matrix_B[188],mul_res1[2588]);
multi_7x28 multi_7x28_mod_2589(clk,rst,matrix_A[2589],matrix_B[189],mul_res1[2589]);
multi_7x28 multi_7x28_mod_2590(clk,rst,matrix_A[2590],matrix_B[190],mul_res1[2590]);
multi_7x28 multi_7x28_mod_2591(clk,rst,matrix_A[2591],matrix_B[191],mul_res1[2591]);
multi_7x28 multi_7x28_mod_2592(clk,rst,matrix_A[2592],matrix_B[192],mul_res1[2592]);
multi_7x28 multi_7x28_mod_2593(clk,rst,matrix_A[2593],matrix_B[193],mul_res1[2593]);
multi_7x28 multi_7x28_mod_2594(clk,rst,matrix_A[2594],matrix_B[194],mul_res1[2594]);
multi_7x28 multi_7x28_mod_2595(clk,rst,matrix_A[2595],matrix_B[195],mul_res1[2595]);
multi_7x28 multi_7x28_mod_2596(clk,rst,matrix_A[2596],matrix_B[196],mul_res1[2596]);
multi_7x28 multi_7x28_mod_2597(clk,rst,matrix_A[2597],matrix_B[197],mul_res1[2597]);
multi_7x28 multi_7x28_mod_2598(clk,rst,matrix_A[2598],matrix_B[198],mul_res1[2598]);
multi_7x28 multi_7x28_mod_2599(clk,rst,matrix_A[2599],matrix_B[199],mul_res1[2599]);
multi_7x28 multi_7x28_mod_2600(clk,rst,matrix_A[2600],matrix_B[0],mul_res1[2600]);
multi_7x28 multi_7x28_mod_2601(clk,rst,matrix_A[2601],matrix_B[1],mul_res1[2601]);
multi_7x28 multi_7x28_mod_2602(clk,rst,matrix_A[2602],matrix_B[2],mul_res1[2602]);
multi_7x28 multi_7x28_mod_2603(clk,rst,matrix_A[2603],matrix_B[3],mul_res1[2603]);
multi_7x28 multi_7x28_mod_2604(clk,rst,matrix_A[2604],matrix_B[4],mul_res1[2604]);
multi_7x28 multi_7x28_mod_2605(clk,rst,matrix_A[2605],matrix_B[5],mul_res1[2605]);
multi_7x28 multi_7x28_mod_2606(clk,rst,matrix_A[2606],matrix_B[6],mul_res1[2606]);
multi_7x28 multi_7x28_mod_2607(clk,rst,matrix_A[2607],matrix_B[7],mul_res1[2607]);
multi_7x28 multi_7x28_mod_2608(clk,rst,matrix_A[2608],matrix_B[8],mul_res1[2608]);
multi_7x28 multi_7x28_mod_2609(clk,rst,matrix_A[2609],matrix_B[9],mul_res1[2609]);
multi_7x28 multi_7x28_mod_2610(clk,rst,matrix_A[2610],matrix_B[10],mul_res1[2610]);
multi_7x28 multi_7x28_mod_2611(clk,rst,matrix_A[2611],matrix_B[11],mul_res1[2611]);
multi_7x28 multi_7x28_mod_2612(clk,rst,matrix_A[2612],matrix_B[12],mul_res1[2612]);
multi_7x28 multi_7x28_mod_2613(clk,rst,matrix_A[2613],matrix_B[13],mul_res1[2613]);
multi_7x28 multi_7x28_mod_2614(clk,rst,matrix_A[2614],matrix_B[14],mul_res1[2614]);
multi_7x28 multi_7x28_mod_2615(clk,rst,matrix_A[2615],matrix_B[15],mul_res1[2615]);
multi_7x28 multi_7x28_mod_2616(clk,rst,matrix_A[2616],matrix_B[16],mul_res1[2616]);
multi_7x28 multi_7x28_mod_2617(clk,rst,matrix_A[2617],matrix_B[17],mul_res1[2617]);
multi_7x28 multi_7x28_mod_2618(clk,rst,matrix_A[2618],matrix_B[18],mul_res1[2618]);
multi_7x28 multi_7x28_mod_2619(clk,rst,matrix_A[2619],matrix_B[19],mul_res1[2619]);
multi_7x28 multi_7x28_mod_2620(clk,rst,matrix_A[2620],matrix_B[20],mul_res1[2620]);
multi_7x28 multi_7x28_mod_2621(clk,rst,matrix_A[2621],matrix_B[21],mul_res1[2621]);
multi_7x28 multi_7x28_mod_2622(clk,rst,matrix_A[2622],matrix_B[22],mul_res1[2622]);
multi_7x28 multi_7x28_mod_2623(clk,rst,matrix_A[2623],matrix_B[23],mul_res1[2623]);
multi_7x28 multi_7x28_mod_2624(clk,rst,matrix_A[2624],matrix_B[24],mul_res1[2624]);
multi_7x28 multi_7x28_mod_2625(clk,rst,matrix_A[2625],matrix_B[25],mul_res1[2625]);
multi_7x28 multi_7x28_mod_2626(clk,rst,matrix_A[2626],matrix_B[26],mul_res1[2626]);
multi_7x28 multi_7x28_mod_2627(clk,rst,matrix_A[2627],matrix_B[27],mul_res1[2627]);
multi_7x28 multi_7x28_mod_2628(clk,rst,matrix_A[2628],matrix_B[28],mul_res1[2628]);
multi_7x28 multi_7x28_mod_2629(clk,rst,matrix_A[2629],matrix_B[29],mul_res1[2629]);
multi_7x28 multi_7x28_mod_2630(clk,rst,matrix_A[2630],matrix_B[30],mul_res1[2630]);
multi_7x28 multi_7x28_mod_2631(clk,rst,matrix_A[2631],matrix_B[31],mul_res1[2631]);
multi_7x28 multi_7x28_mod_2632(clk,rst,matrix_A[2632],matrix_B[32],mul_res1[2632]);
multi_7x28 multi_7x28_mod_2633(clk,rst,matrix_A[2633],matrix_B[33],mul_res1[2633]);
multi_7x28 multi_7x28_mod_2634(clk,rst,matrix_A[2634],matrix_B[34],mul_res1[2634]);
multi_7x28 multi_7x28_mod_2635(clk,rst,matrix_A[2635],matrix_B[35],mul_res1[2635]);
multi_7x28 multi_7x28_mod_2636(clk,rst,matrix_A[2636],matrix_B[36],mul_res1[2636]);
multi_7x28 multi_7x28_mod_2637(clk,rst,matrix_A[2637],matrix_B[37],mul_res1[2637]);
multi_7x28 multi_7x28_mod_2638(clk,rst,matrix_A[2638],matrix_B[38],mul_res1[2638]);
multi_7x28 multi_7x28_mod_2639(clk,rst,matrix_A[2639],matrix_B[39],mul_res1[2639]);
multi_7x28 multi_7x28_mod_2640(clk,rst,matrix_A[2640],matrix_B[40],mul_res1[2640]);
multi_7x28 multi_7x28_mod_2641(clk,rst,matrix_A[2641],matrix_B[41],mul_res1[2641]);
multi_7x28 multi_7x28_mod_2642(clk,rst,matrix_A[2642],matrix_B[42],mul_res1[2642]);
multi_7x28 multi_7x28_mod_2643(clk,rst,matrix_A[2643],matrix_B[43],mul_res1[2643]);
multi_7x28 multi_7x28_mod_2644(clk,rst,matrix_A[2644],matrix_B[44],mul_res1[2644]);
multi_7x28 multi_7x28_mod_2645(clk,rst,matrix_A[2645],matrix_B[45],mul_res1[2645]);
multi_7x28 multi_7x28_mod_2646(clk,rst,matrix_A[2646],matrix_B[46],mul_res1[2646]);
multi_7x28 multi_7x28_mod_2647(clk,rst,matrix_A[2647],matrix_B[47],mul_res1[2647]);
multi_7x28 multi_7x28_mod_2648(clk,rst,matrix_A[2648],matrix_B[48],mul_res1[2648]);
multi_7x28 multi_7x28_mod_2649(clk,rst,matrix_A[2649],matrix_B[49],mul_res1[2649]);
multi_7x28 multi_7x28_mod_2650(clk,rst,matrix_A[2650],matrix_B[50],mul_res1[2650]);
multi_7x28 multi_7x28_mod_2651(clk,rst,matrix_A[2651],matrix_B[51],mul_res1[2651]);
multi_7x28 multi_7x28_mod_2652(clk,rst,matrix_A[2652],matrix_B[52],mul_res1[2652]);
multi_7x28 multi_7x28_mod_2653(clk,rst,matrix_A[2653],matrix_B[53],mul_res1[2653]);
multi_7x28 multi_7x28_mod_2654(clk,rst,matrix_A[2654],matrix_B[54],mul_res1[2654]);
multi_7x28 multi_7x28_mod_2655(clk,rst,matrix_A[2655],matrix_B[55],mul_res1[2655]);
multi_7x28 multi_7x28_mod_2656(clk,rst,matrix_A[2656],matrix_B[56],mul_res1[2656]);
multi_7x28 multi_7x28_mod_2657(clk,rst,matrix_A[2657],matrix_B[57],mul_res1[2657]);
multi_7x28 multi_7x28_mod_2658(clk,rst,matrix_A[2658],matrix_B[58],mul_res1[2658]);
multi_7x28 multi_7x28_mod_2659(clk,rst,matrix_A[2659],matrix_B[59],mul_res1[2659]);
multi_7x28 multi_7x28_mod_2660(clk,rst,matrix_A[2660],matrix_B[60],mul_res1[2660]);
multi_7x28 multi_7x28_mod_2661(clk,rst,matrix_A[2661],matrix_B[61],mul_res1[2661]);
multi_7x28 multi_7x28_mod_2662(clk,rst,matrix_A[2662],matrix_B[62],mul_res1[2662]);
multi_7x28 multi_7x28_mod_2663(clk,rst,matrix_A[2663],matrix_B[63],mul_res1[2663]);
multi_7x28 multi_7x28_mod_2664(clk,rst,matrix_A[2664],matrix_B[64],mul_res1[2664]);
multi_7x28 multi_7x28_mod_2665(clk,rst,matrix_A[2665],matrix_B[65],mul_res1[2665]);
multi_7x28 multi_7x28_mod_2666(clk,rst,matrix_A[2666],matrix_B[66],mul_res1[2666]);
multi_7x28 multi_7x28_mod_2667(clk,rst,matrix_A[2667],matrix_B[67],mul_res1[2667]);
multi_7x28 multi_7x28_mod_2668(clk,rst,matrix_A[2668],matrix_B[68],mul_res1[2668]);
multi_7x28 multi_7x28_mod_2669(clk,rst,matrix_A[2669],matrix_B[69],mul_res1[2669]);
multi_7x28 multi_7x28_mod_2670(clk,rst,matrix_A[2670],matrix_B[70],mul_res1[2670]);
multi_7x28 multi_7x28_mod_2671(clk,rst,matrix_A[2671],matrix_B[71],mul_res1[2671]);
multi_7x28 multi_7x28_mod_2672(clk,rst,matrix_A[2672],matrix_B[72],mul_res1[2672]);
multi_7x28 multi_7x28_mod_2673(clk,rst,matrix_A[2673],matrix_B[73],mul_res1[2673]);
multi_7x28 multi_7x28_mod_2674(clk,rst,matrix_A[2674],matrix_B[74],mul_res1[2674]);
multi_7x28 multi_7x28_mod_2675(clk,rst,matrix_A[2675],matrix_B[75],mul_res1[2675]);
multi_7x28 multi_7x28_mod_2676(clk,rst,matrix_A[2676],matrix_B[76],mul_res1[2676]);
multi_7x28 multi_7x28_mod_2677(clk,rst,matrix_A[2677],matrix_B[77],mul_res1[2677]);
multi_7x28 multi_7x28_mod_2678(clk,rst,matrix_A[2678],matrix_B[78],mul_res1[2678]);
multi_7x28 multi_7x28_mod_2679(clk,rst,matrix_A[2679],matrix_B[79],mul_res1[2679]);
multi_7x28 multi_7x28_mod_2680(clk,rst,matrix_A[2680],matrix_B[80],mul_res1[2680]);
multi_7x28 multi_7x28_mod_2681(clk,rst,matrix_A[2681],matrix_B[81],mul_res1[2681]);
multi_7x28 multi_7x28_mod_2682(clk,rst,matrix_A[2682],matrix_B[82],mul_res1[2682]);
multi_7x28 multi_7x28_mod_2683(clk,rst,matrix_A[2683],matrix_B[83],mul_res1[2683]);
multi_7x28 multi_7x28_mod_2684(clk,rst,matrix_A[2684],matrix_B[84],mul_res1[2684]);
multi_7x28 multi_7x28_mod_2685(clk,rst,matrix_A[2685],matrix_B[85],mul_res1[2685]);
multi_7x28 multi_7x28_mod_2686(clk,rst,matrix_A[2686],matrix_B[86],mul_res1[2686]);
multi_7x28 multi_7x28_mod_2687(clk,rst,matrix_A[2687],matrix_B[87],mul_res1[2687]);
multi_7x28 multi_7x28_mod_2688(clk,rst,matrix_A[2688],matrix_B[88],mul_res1[2688]);
multi_7x28 multi_7x28_mod_2689(clk,rst,matrix_A[2689],matrix_B[89],mul_res1[2689]);
multi_7x28 multi_7x28_mod_2690(clk,rst,matrix_A[2690],matrix_B[90],mul_res1[2690]);
multi_7x28 multi_7x28_mod_2691(clk,rst,matrix_A[2691],matrix_B[91],mul_res1[2691]);
multi_7x28 multi_7x28_mod_2692(clk,rst,matrix_A[2692],matrix_B[92],mul_res1[2692]);
multi_7x28 multi_7x28_mod_2693(clk,rst,matrix_A[2693],matrix_B[93],mul_res1[2693]);
multi_7x28 multi_7x28_mod_2694(clk,rst,matrix_A[2694],matrix_B[94],mul_res1[2694]);
multi_7x28 multi_7x28_mod_2695(clk,rst,matrix_A[2695],matrix_B[95],mul_res1[2695]);
multi_7x28 multi_7x28_mod_2696(clk,rst,matrix_A[2696],matrix_B[96],mul_res1[2696]);
multi_7x28 multi_7x28_mod_2697(clk,rst,matrix_A[2697],matrix_B[97],mul_res1[2697]);
multi_7x28 multi_7x28_mod_2698(clk,rst,matrix_A[2698],matrix_B[98],mul_res1[2698]);
multi_7x28 multi_7x28_mod_2699(clk,rst,matrix_A[2699],matrix_B[99],mul_res1[2699]);
multi_7x28 multi_7x28_mod_2700(clk,rst,matrix_A[2700],matrix_B[100],mul_res1[2700]);
multi_7x28 multi_7x28_mod_2701(clk,rst,matrix_A[2701],matrix_B[101],mul_res1[2701]);
multi_7x28 multi_7x28_mod_2702(clk,rst,matrix_A[2702],matrix_B[102],mul_res1[2702]);
multi_7x28 multi_7x28_mod_2703(clk,rst,matrix_A[2703],matrix_B[103],mul_res1[2703]);
multi_7x28 multi_7x28_mod_2704(clk,rst,matrix_A[2704],matrix_B[104],mul_res1[2704]);
multi_7x28 multi_7x28_mod_2705(clk,rst,matrix_A[2705],matrix_B[105],mul_res1[2705]);
multi_7x28 multi_7x28_mod_2706(clk,rst,matrix_A[2706],matrix_B[106],mul_res1[2706]);
multi_7x28 multi_7x28_mod_2707(clk,rst,matrix_A[2707],matrix_B[107],mul_res1[2707]);
multi_7x28 multi_7x28_mod_2708(clk,rst,matrix_A[2708],matrix_B[108],mul_res1[2708]);
multi_7x28 multi_7x28_mod_2709(clk,rst,matrix_A[2709],matrix_B[109],mul_res1[2709]);
multi_7x28 multi_7x28_mod_2710(clk,rst,matrix_A[2710],matrix_B[110],mul_res1[2710]);
multi_7x28 multi_7x28_mod_2711(clk,rst,matrix_A[2711],matrix_B[111],mul_res1[2711]);
multi_7x28 multi_7x28_mod_2712(clk,rst,matrix_A[2712],matrix_B[112],mul_res1[2712]);
multi_7x28 multi_7x28_mod_2713(clk,rst,matrix_A[2713],matrix_B[113],mul_res1[2713]);
multi_7x28 multi_7x28_mod_2714(clk,rst,matrix_A[2714],matrix_B[114],mul_res1[2714]);
multi_7x28 multi_7x28_mod_2715(clk,rst,matrix_A[2715],matrix_B[115],mul_res1[2715]);
multi_7x28 multi_7x28_mod_2716(clk,rst,matrix_A[2716],matrix_B[116],mul_res1[2716]);
multi_7x28 multi_7x28_mod_2717(clk,rst,matrix_A[2717],matrix_B[117],mul_res1[2717]);
multi_7x28 multi_7x28_mod_2718(clk,rst,matrix_A[2718],matrix_B[118],mul_res1[2718]);
multi_7x28 multi_7x28_mod_2719(clk,rst,matrix_A[2719],matrix_B[119],mul_res1[2719]);
multi_7x28 multi_7x28_mod_2720(clk,rst,matrix_A[2720],matrix_B[120],mul_res1[2720]);
multi_7x28 multi_7x28_mod_2721(clk,rst,matrix_A[2721],matrix_B[121],mul_res1[2721]);
multi_7x28 multi_7x28_mod_2722(clk,rst,matrix_A[2722],matrix_B[122],mul_res1[2722]);
multi_7x28 multi_7x28_mod_2723(clk,rst,matrix_A[2723],matrix_B[123],mul_res1[2723]);
multi_7x28 multi_7x28_mod_2724(clk,rst,matrix_A[2724],matrix_B[124],mul_res1[2724]);
multi_7x28 multi_7x28_mod_2725(clk,rst,matrix_A[2725],matrix_B[125],mul_res1[2725]);
multi_7x28 multi_7x28_mod_2726(clk,rst,matrix_A[2726],matrix_B[126],mul_res1[2726]);
multi_7x28 multi_7x28_mod_2727(clk,rst,matrix_A[2727],matrix_B[127],mul_res1[2727]);
multi_7x28 multi_7x28_mod_2728(clk,rst,matrix_A[2728],matrix_B[128],mul_res1[2728]);
multi_7x28 multi_7x28_mod_2729(clk,rst,matrix_A[2729],matrix_B[129],mul_res1[2729]);
multi_7x28 multi_7x28_mod_2730(clk,rst,matrix_A[2730],matrix_B[130],mul_res1[2730]);
multi_7x28 multi_7x28_mod_2731(clk,rst,matrix_A[2731],matrix_B[131],mul_res1[2731]);
multi_7x28 multi_7x28_mod_2732(clk,rst,matrix_A[2732],matrix_B[132],mul_res1[2732]);
multi_7x28 multi_7x28_mod_2733(clk,rst,matrix_A[2733],matrix_B[133],mul_res1[2733]);
multi_7x28 multi_7x28_mod_2734(clk,rst,matrix_A[2734],matrix_B[134],mul_res1[2734]);
multi_7x28 multi_7x28_mod_2735(clk,rst,matrix_A[2735],matrix_B[135],mul_res1[2735]);
multi_7x28 multi_7x28_mod_2736(clk,rst,matrix_A[2736],matrix_B[136],mul_res1[2736]);
multi_7x28 multi_7x28_mod_2737(clk,rst,matrix_A[2737],matrix_B[137],mul_res1[2737]);
multi_7x28 multi_7x28_mod_2738(clk,rst,matrix_A[2738],matrix_B[138],mul_res1[2738]);
multi_7x28 multi_7x28_mod_2739(clk,rst,matrix_A[2739],matrix_B[139],mul_res1[2739]);
multi_7x28 multi_7x28_mod_2740(clk,rst,matrix_A[2740],matrix_B[140],mul_res1[2740]);
multi_7x28 multi_7x28_mod_2741(clk,rst,matrix_A[2741],matrix_B[141],mul_res1[2741]);
multi_7x28 multi_7x28_mod_2742(clk,rst,matrix_A[2742],matrix_B[142],mul_res1[2742]);
multi_7x28 multi_7x28_mod_2743(clk,rst,matrix_A[2743],matrix_B[143],mul_res1[2743]);
multi_7x28 multi_7x28_mod_2744(clk,rst,matrix_A[2744],matrix_B[144],mul_res1[2744]);
multi_7x28 multi_7x28_mod_2745(clk,rst,matrix_A[2745],matrix_B[145],mul_res1[2745]);
multi_7x28 multi_7x28_mod_2746(clk,rst,matrix_A[2746],matrix_B[146],mul_res1[2746]);
multi_7x28 multi_7x28_mod_2747(clk,rst,matrix_A[2747],matrix_B[147],mul_res1[2747]);
multi_7x28 multi_7x28_mod_2748(clk,rst,matrix_A[2748],matrix_B[148],mul_res1[2748]);
multi_7x28 multi_7x28_mod_2749(clk,rst,matrix_A[2749],matrix_B[149],mul_res1[2749]);
multi_7x28 multi_7x28_mod_2750(clk,rst,matrix_A[2750],matrix_B[150],mul_res1[2750]);
multi_7x28 multi_7x28_mod_2751(clk,rst,matrix_A[2751],matrix_B[151],mul_res1[2751]);
multi_7x28 multi_7x28_mod_2752(clk,rst,matrix_A[2752],matrix_B[152],mul_res1[2752]);
multi_7x28 multi_7x28_mod_2753(clk,rst,matrix_A[2753],matrix_B[153],mul_res1[2753]);
multi_7x28 multi_7x28_mod_2754(clk,rst,matrix_A[2754],matrix_B[154],mul_res1[2754]);
multi_7x28 multi_7x28_mod_2755(clk,rst,matrix_A[2755],matrix_B[155],mul_res1[2755]);
multi_7x28 multi_7x28_mod_2756(clk,rst,matrix_A[2756],matrix_B[156],mul_res1[2756]);
multi_7x28 multi_7x28_mod_2757(clk,rst,matrix_A[2757],matrix_B[157],mul_res1[2757]);
multi_7x28 multi_7x28_mod_2758(clk,rst,matrix_A[2758],matrix_B[158],mul_res1[2758]);
multi_7x28 multi_7x28_mod_2759(clk,rst,matrix_A[2759],matrix_B[159],mul_res1[2759]);
multi_7x28 multi_7x28_mod_2760(clk,rst,matrix_A[2760],matrix_B[160],mul_res1[2760]);
multi_7x28 multi_7x28_mod_2761(clk,rst,matrix_A[2761],matrix_B[161],mul_res1[2761]);
multi_7x28 multi_7x28_mod_2762(clk,rst,matrix_A[2762],matrix_B[162],mul_res1[2762]);
multi_7x28 multi_7x28_mod_2763(clk,rst,matrix_A[2763],matrix_B[163],mul_res1[2763]);
multi_7x28 multi_7x28_mod_2764(clk,rst,matrix_A[2764],matrix_B[164],mul_res1[2764]);
multi_7x28 multi_7x28_mod_2765(clk,rst,matrix_A[2765],matrix_B[165],mul_res1[2765]);
multi_7x28 multi_7x28_mod_2766(clk,rst,matrix_A[2766],matrix_B[166],mul_res1[2766]);
multi_7x28 multi_7x28_mod_2767(clk,rst,matrix_A[2767],matrix_B[167],mul_res1[2767]);
multi_7x28 multi_7x28_mod_2768(clk,rst,matrix_A[2768],matrix_B[168],mul_res1[2768]);
multi_7x28 multi_7x28_mod_2769(clk,rst,matrix_A[2769],matrix_B[169],mul_res1[2769]);
multi_7x28 multi_7x28_mod_2770(clk,rst,matrix_A[2770],matrix_B[170],mul_res1[2770]);
multi_7x28 multi_7x28_mod_2771(clk,rst,matrix_A[2771],matrix_B[171],mul_res1[2771]);
multi_7x28 multi_7x28_mod_2772(clk,rst,matrix_A[2772],matrix_B[172],mul_res1[2772]);
multi_7x28 multi_7x28_mod_2773(clk,rst,matrix_A[2773],matrix_B[173],mul_res1[2773]);
multi_7x28 multi_7x28_mod_2774(clk,rst,matrix_A[2774],matrix_B[174],mul_res1[2774]);
multi_7x28 multi_7x28_mod_2775(clk,rst,matrix_A[2775],matrix_B[175],mul_res1[2775]);
multi_7x28 multi_7x28_mod_2776(clk,rst,matrix_A[2776],matrix_B[176],mul_res1[2776]);
multi_7x28 multi_7x28_mod_2777(clk,rst,matrix_A[2777],matrix_B[177],mul_res1[2777]);
multi_7x28 multi_7x28_mod_2778(clk,rst,matrix_A[2778],matrix_B[178],mul_res1[2778]);
multi_7x28 multi_7x28_mod_2779(clk,rst,matrix_A[2779],matrix_B[179],mul_res1[2779]);
multi_7x28 multi_7x28_mod_2780(clk,rst,matrix_A[2780],matrix_B[180],mul_res1[2780]);
multi_7x28 multi_7x28_mod_2781(clk,rst,matrix_A[2781],matrix_B[181],mul_res1[2781]);
multi_7x28 multi_7x28_mod_2782(clk,rst,matrix_A[2782],matrix_B[182],mul_res1[2782]);
multi_7x28 multi_7x28_mod_2783(clk,rst,matrix_A[2783],matrix_B[183],mul_res1[2783]);
multi_7x28 multi_7x28_mod_2784(clk,rst,matrix_A[2784],matrix_B[184],mul_res1[2784]);
multi_7x28 multi_7x28_mod_2785(clk,rst,matrix_A[2785],matrix_B[185],mul_res1[2785]);
multi_7x28 multi_7x28_mod_2786(clk,rst,matrix_A[2786],matrix_B[186],mul_res1[2786]);
multi_7x28 multi_7x28_mod_2787(clk,rst,matrix_A[2787],matrix_B[187],mul_res1[2787]);
multi_7x28 multi_7x28_mod_2788(clk,rst,matrix_A[2788],matrix_B[188],mul_res1[2788]);
multi_7x28 multi_7x28_mod_2789(clk,rst,matrix_A[2789],matrix_B[189],mul_res1[2789]);
multi_7x28 multi_7x28_mod_2790(clk,rst,matrix_A[2790],matrix_B[190],mul_res1[2790]);
multi_7x28 multi_7x28_mod_2791(clk,rst,matrix_A[2791],matrix_B[191],mul_res1[2791]);
multi_7x28 multi_7x28_mod_2792(clk,rst,matrix_A[2792],matrix_B[192],mul_res1[2792]);
multi_7x28 multi_7x28_mod_2793(clk,rst,matrix_A[2793],matrix_B[193],mul_res1[2793]);
multi_7x28 multi_7x28_mod_2794(clk,rst,matrix_A[2794],matrix_B[194],mul_res1[2794]);
multi_7x28 multi_7x28_mod_2795(clk,rst,matrix_A[2795],matrix_B[195],mul_res1[2795]);
multi_7x28 multi_7x28_mod_2796(clk,rst,matrix_A[2796],matrix_B[196],mul_res1[2796]);
multi_7x28 multi_7x28_mod_2797(clk,rst,matrix_A[2797],matrix_B[197],mul_res1[2797]);
multi_7x28 multi_7x28_mod_2798(clk,rst,matrix_A[2798],matrix_B[198],mul_res1[2798]);
multi_7x28 multi_7x28_mod_2799(clk,rst,matrix_A[2799],matrix_B[199],mul_res1[2799]);
multi_7x28 multi_7x28_mod_2800(clk,rst,matrix_A[2800],matrix_B[0],mul_res1[2800]);
multi_7x28 multi_7x28_mod_2801(clk,rst,matrix_A[2801],matrix_B[1],mul_res1[2801]);
multi_7x28 multi_7x28_mod_2802(clk,rst,matrix_A[2802],matrix_B[2],mul_res1[2802]);
multi_7x28 multi_7x28_mod_2803(clk,rst,matrix_A[2803],matrix_B[3],mul_res1[2803]);
multi_7x28 multi_7x28_mod_2804(clk,rst,matrix_A[2804],matrix_B[4],mul_res1[2804]);
multi_7x28 multi_7x28_mod_2805(clk,rst,matrix_A[2805],matrix_B[5],mul_res1[2805]);
multi_7x28 multi_7x28_mod_2806(clk,rst,matrix_A[2806],matrix_B[6],mul_res1[2806]);
multi_7x28 multi_7x28_mod_2807(clk,rst,matrix_A[2807],matrix_B[7],mul_res1[2807]);
multi_7x28 multi_7x28_mod_2808(clk,rst,matrix_A[2808],matrix_B[8],mul_res1[2808]);
multi_7x28 multi_7x28_mod_2809(clk,rst,matrix_A[2809],matrix_B[9],mul_res1[2809]);
multi_7x28 multi_7x28_mod_2810(clk,rst,matrix_A[2810],matrix_B[10],mul_res1[2810]);
multi_7x28 multi_7x28_mod_2811(clk,rst,matrix_A[2811],matrix_B[11],mul_res1[2811]);
multi_7x28 multi_7x28_mod_2812(clk,rst,matrix_A[2812],matrix_B[12],mul_res1[2812]);
multi_7x28 multi_7x28_mod_2813(clk,rst,matrix_A[2813],matrix_B[13],mul_res1[2813]);
multi_7x28 multi_7x28_mod_2814(clk,rst,matrix_A[2814],matrix_B[14],mul_res1[2814]);
multi_7x28 multi_7x28_mod_2815(clk,rst,matrix_A[2815],matrix_B[15],mul_res1[2815]);
multi_7x28 multi_7x28_mod_2816(clk,rst,matrix_A[2816],matrix_B[16],mul_res1[2816]);
multi_7x28 multi_7x28_mod_2817(clk,rst,matrix_A[2817],matrix_B[17],mul_res1[2817]);
multi_7x28 multi_7x28_mod_2818(clk,rst,matrix_A[2818],matrix_B[18],mul_res1[2818]);
multi_7x28 multi_7x28_mod_2819(clk,rst,matrix_A[2819],matrix_B[19],mul_res1[2819]);
multi_7x28 multi_7x28_mod_2820(clk,rst,matrix_A[2820],matrix_B[20],mul_res1[2820]);
multi_7x28 multi_7x28_mod_2821(clk,rst,matrix_A[2821],matrix_B[21],mul_res1[2821]);
multi_7x28 multi_7x28_mod_2822(clk,rst,matrix_A[2822],matrix_B[22],mul_res1[2822]);
multi_7x28 multi_7x28_mod_2823(clk,rst,matrix_A[2823],matrix_B[23],mul_res1[2823]);
multi_7x28 multi_7x28_mod_2824(clk,rst,matrix_A[2824],matrix_B[24],mul_res1[2824]);
multi_7x28 multi_7x28_mod_2825(clk,rst,matrix_A[2825],matrix_B[25],mul_res1[2825]);
multi_7x28 multi_7x28_mod_2826(clk,rst,matrix_A[2826],matrix_B[26],mul_res1[2826]);
multi_7x28 multi_7x28_mod_2827(clk,rst,matrix_A[2827],matrix_B[27],mul_res1[2827]);
multi_7x28 multi_7x28_mod_2828(clk,rst,matrix_A[2828],matrix_B[28],mul_res1[2828]);
multi_7x28 multi_7x28_mod_2829(clk,rst,matrix_A[2829],matrix_B[29],mul_res1[2829]);
multi_7x28 multi_7x28_mod_2830(clk,rst,matrix_A[2830],matrix_B[30],mul_res1[2830]);
multi_7x28 multi_7x28_mod_2831(clk,rst,matrix_A[2831],matrix_B[31],mul_res1[2831]);
multi_7x28 multi_7x28_mod_2832(clk,rst,matrix_A[2832],matrix_B[32],mul_res1[2832]);
multi_7x28 multi_7x28_mod_2833(clk,rst,matrix_A[2833],matrix_B[33],mul_res1[2833]);
multi_7x28 multi_7x28_mod_2834(clk,rst,matrix_A[2834],matrix_B[34],mul_res1[2834]);
multi_7x28 multi_7x28_mod_2835(clk,rst,matrix_A[2835],matrix_B[35],mul_res1[2835]);
multi_7x28 multi_7x28_mod_2836(clk,rst,matrix_A[2836],matrix_B[36],mul_res1[2836]);
multi_7x28 multi_7x28_mod_2837(clk,rst,matrix_A[2837],matrix_B[37],mul_res1[2837]);
multi_7x28 multi_7x28_mod_2838(clk,rst,matrix_A[2838],matrix_B[38],mul_res1[2838]);
multi_7x28 multi_7x28_mod_2839(clk,rst,matrix_A[2839],matrix_B[39],mul_res1[2839]);
multi_7x28 multi_7x28_mod_2840(clk,rst,matrix_A[2840],matrix_B[40],mul_res1[2840]);
multi_7x28 multi_7x28_mod_2841(clk,rst,matrix_A[2841],matrix_B[41],mul_res1[2841]);
multi_7x28 multi_7x28_mod_2842(clk,rst,matrix_A[2842],matrix_B[42],mul_res1[2842]);
multi_7x28 multi_7x28_mod_2843(clk,rst,matrix_A[2843],matrix_B[43],mul_res1[2843]);
multi_7x28 multi_7x28_mod_2844(clk,rst,matrix_A[2844],matrix_B[44],mul_res1[2844]);
multi_7x28 multi_7x28_mod_2845(clk,rst,matrix_A[2845],matrix_B[45],mul_res1[2845]);
multi_7x28 multi_7x28_mod_2846(clk,rst,matrix_A[2846],matrix_B[46],mul_res1[2846]);
multi_7x28 multi_7x28_mod_2847(clk,rst,matrix_A[2847],matrix_B[47],mul_res1[2847]);
multi_7x28 multi_7x28_mod_2848(clk,rst,matrix_A[2848],matrix_B[48],mul_res1[2848]);
multi_7x28 multi_7x28_mod_2849(clk,rst,matrix_A[2849],matrix_B[49],mul_res1[2849]);
multi_7x28 multi_7x28_mod_2850(clk,rst,matrix_A[2850],matrix_B[50],mul_res1[2850]);
multi_7x28 multi_7x28_mod_2851(clk,rst,matrix_A[2851],matrix_B[51],mul_res1[2851]);
multi_7x28 multi_7x28_mod_2852(clk,rst,matrix_A[2852],matrix_B[52],mul_res1[2852]);
multi_7x28 multi_7x28_mod_2853(clk,rst,matrix_A[2853],matrix_B[53],mul_res1[2853]);
multi_7x28 multi_7x28_mod_2854(clk,rst,matrix_A[2854],matrix_B[54],mul_res1[2854]);
multi_7x28 multi_7x28_mod_2855(clk,rst,matrix_A[2855],matrix_B[55],mul_res1[2855]);
multi_7x28 multi_7x28_mod_2856(clk,rst,matrix_A[2856],matrix_B[56],mul_res1[2856]);
multi_7x28 multi_7x28_mod_2857(clk,rst,matrix_A[2857],matrix_B[57],mul_res1[2857]);
multi_7x28 multi_7x28_mod_2858(clk,rst,matrix_A[2858],matrix_B[58],mul_res1[2858]);
multi_7x28 multi_7x28_mod_2859(clk,rst,matrix_A[2859],matrix_B[59],mul_res1[2859]);
multi_7x28 multi_7x28_mod_2860(clk,rst,matrix_A[2860],matrix_B[60],mul_res1[2860]);
multi_7x28 multi_7x28_mod_2861(clk,rst,matrix_A[2861],matrix_B[61],mul_res1[2861]);
multi_7x28 multi_7x28_mod_2862(clk,rst,matrix_A[2862],matrix_B[62],mul_res1[2862]);
multi_7x28 multi_7x28_mod_2863(clk,rst,matrix_A[2863],matrix_B[63],mul_res1[2863]);
multi_7x28 multi_7x28_mod_2864(clk,rst,matrix_A[2864],matrix_B[64],mul_res1[2864]);
multi_7x28 multi_7x28_mod_2865(clk,rst,matrix_A[2865],matrix_B[65],mul_res1[2865]);
multi_7x28 multi_7x28_mod_2866(clk,rst,matrix_A[2866],matrix_B[66],mul_res1[2866]);
multi_7x28 multi_7x28_mod_2867(clk,rst,matrix_A[2867],matrix_B[67],mul_res1[2867]);
multi_7x28 multi_7x28_mod_2868(clk,rst,matrix_A[2868],matrix_B[68],mul_res1[2868]);
multi_7x28 multi_7x28_mod_2869(clk,rst,matrix_A[2869],matrix_B[69],mul_res1[2869]);
multi_7x28 multi_7x28_mod_2870(clk,rst,matrix_A[2870],matrix_B[70],mul_res1[2870]);
multi_7x28 multi_7x28_mod_2871(clk,rst,matrix_A[2871],matrix_B[71],mul_res1[2871]);
multi_7x28 multi_7x28_mod_2872(clk,rst,matrix_A[2872],matrix_B[72],mul_res1[2872]);
multi_7x28 multi_7x28_mod_2873(clk,rst,matrix_A[2873],matrix_B[73],mul_res1[2873]);
multi_7x28 multi_7x28_mod_2874(clk,rst,matrix_A[2874],matrix_B[74],mul_res1[2874]);
multi_7x28 multi_7x28_mod_2875(clk,rst,matrix_A[2875],matrix_B[75],mul_res1[2875]);
multi_7x28 multi_7x28_mod_2876(clk,rst,matrix_A[2876],matrix_B[76],mul_res1[2876]);
multi_7x28 multi_7x28_mod_2877(clk,rst,matrix_A[2877],matrix_B[77],mul_res1[2877]);
multi_7x28 multi_7x28_mod_2878(clk,rst,matrix_A[2878],matrix_B[78],mul_res1[2878]);
multi_7x28 multi_7x28_mod_2879(clk,rst,matrix_A[2879],matrix_B[79],mul_res1[2879]);
multi_7x28 multi_7x28_mod_2880(clk,rst,matrix_A[2880],matrix_B[80],mul_res1[2880]);
multi_7x28 multi_7x28_mod_2881(clk,rst,matrix_A[2881],matrix_B[81],mul_res1[2881]);
multi_7x28 multi_7x28_mod_2882(clk,rst,matrix_A[2882],matrix_B[82],mul_res1[2882]);
multi_7x28 multi_7x28_mod_2883(clk,rst,matrix_A[2883],matrix_B[83],mul_res1[2883]);
multi_7x28 multi_7x28_mod_2884(clk,rst,matrix_A[2884],matrix_B[84],mul_res1[2884]);
multi_7x28 multi_7x28_mod_2885(clk,rst,matrix_A[2885],matrix_B[85],mul_res1[2885]);
multi_7x28 multi_7x28_mod_2886(clk,rst,matrix_A[2886],matrix_B[86],mul_res1[2886]);
multi_7x28 multi_7x28_mod_2887(clk,rst,matrix_A[2887],matrix_B[87],mul_res1[2887]);
multi_7x28 multi_7x28_mod_2888(clk,rst,matrix_A[2888],matrix_B[88],mul_res1[2888]);
multi_7x28 multi_7x28_mod_2889(clk,rst,matrix_A[2889],matrix_B[89],mul_res1[2889]);
multi_7x28 multi_7x28_mod_2890(clk,rst,matrix_A[2890],matrix_B[90],mul_res1[2890]);
multi_7x28 multi_7x28_mod_2891(clk,rst,matrix_A[2891],matrix_B[91],mul_res1[2891]);
multi_7x28 multi_7x28_mod_2892(clk,rst,matrix_A[2892],matrix_B[92],mul_res1[2892]);
multi_7x28 multi_7x28_mod_2893(clk,rst,matrix_A[2893],matrix_B[93],mul_res1[2893]);
multi_7x28 multi_7x28_mod_2894(clk,rst,matrix_A[2894],matrix_B[94],mul_res1[2894]);
multi_7x28 multi_7x28_mod_2895(clk,rst,matrix_A[2895],matrix_B[95],mul_res1[2895]);
multi_7x28 multi_7x28_mod_2896(clk,rst,matrix_A[2896],matrix_B[96],mul_res1[2896]);
multi_7x28 multi_7x28_mod_2897(clk,rst,matrix_A[2897],matrix_B[97],mul_res1[2897]);
multi_7x28 multi_7x28_mod_2898(clk,rst,matrix_A[2898],matrix_B[98],mul_res1[2898]);
multi_7x28 multi_7x28_mod_2899(clk,rst,matrix_A[2899],matrix_B[99],mul_res1[2899]);
multi_7x28 multi_7x28_mod_2900(clk,rst,matrix_A[2900],matrix_B[100],mul_res1[2900]);
multi_7x28 multi_7x28_mod_2901(clk,rst,matrix_A[2901],matrix_B[101],mul_res1[2901]);
multi_7x28 multi_7x28_mod_2902(clk,rst,matrix_A[2902],matrix_B[102],mul_res1[2902]);
multi_7x28 multi_7x28_mod_2903(clk,rst,matrix_A[2903],matrix_B[103],mul_res1[2903]);
multi_7x28 multi_7x28_mod_2904(clk,rst,matrix_A[2904],matrix_B[104],mul_res1[2904]);
multi_7x28 multi_7x28_mod_2905(clk,rst,matrix_A[2905],matrix_B[105],mul_res1[2905]);
multi_7x28 multi_7x28_mod_2906(clk,rst,matrix_A[2906],matrix_B[106],mul_res1[2906]);
multi_7x28 multi_7x28_mod_2907(clk,rst,matrix_A[2907],matrix_B[107],mul_res1[2907]);
multi_7x28 multi_7x28_mod_2908(clk,rst,matrix_A[2908],matrix_B[108],mul_res1[2908]);
multi_7x28 multi_7x28_mod_2909(clk,rst,matrix_A[2909],matrix_B[109],mul_res1[2909]);
multi_7x28 multi_7x28_mod_2910(clk,rst,matrix_A[2910],matrix_B[110],mul_res1[2910]);
multi_7x28 multi_7x28_mod_2911(clk,rst,matrix_A[2911],matrix_B[111],mul_res1[2911]);
multi_7x28 multi_7x28_mod_2912(clk,rst,matrix_A[2912],matrix_B[112],mul_res1[2912]);
multi_7x28 multi_7x28_mod_2913(clk,rst,matrix_A[2913],matrix_B[113],mul_res1[2913]);
multi_7x28 multi_7x28_mod_2914(clk,rst,matrix_A[2914],matrix_B[114],mul_res1[2914]);
multi_7x28 multi_7x28_mod_2915(clk,rst,matrix_A[2915],matrix_B[115],mul_res1[2915]);
multi_7x28 multi_7x28_mod_2916(clk,rst,matrix_A[2916],matrix_B[116],mul_res1[2916]);
multi_7x28 multi_7x28_mod_2917(clk,rst,matrix_A[2917],matrix_B[117],mul_res1[2917]);
multi_7x28 multi_7x28_mod_2918(clk,rst,matrix_A[2918],matrix_B[118],mul_res1[2918]);
multi_7x28 multi_7x28_mod_2919(clk,rst,matrix_A[2919],matrix_B[119],mul_res1[2919]);
multi_7x28 multi_7x28_mod_2920(clk,rst,matrix_A[2920],matrix_B[120],mul_res1[2920]);
multi_7x28 multi_7x28_mod_2921(clk,rst,matrix_A[2921],matrix_B[121],mul_res1[2921]);
multi_7x28 multi_7x28_mod_2922(clk,rst,matrix_A[2922],matrix_B[122],mul_res1[2922]);
multi_7x28 multi_7x28_mod_2923(clk,rst,matrix_A[2923],matrix_B[123],mul_res1[2923]);
multi_7x28 multi_7x28_mod_2924(clk,rst,matrix_A[2924],matrix_B[124],mul_res1[2924]);
multi_7x28 multi_7x28_mod_2925(clk,rst,matrix_A[2925],matrix_B[125],mul_res1[2925]);
multi_7x28 multi_7x28_mod_2926(clk,rst,matrix_A[2926],matrix_B[126],mul_res1[2926]);
multi_7x28 multi_7x28_mod_2927(clk,rst,matrix_A[2927],matrix_B[127],mul_res1[2927]);
multi_7x28 multi_7x28_mod_2928(clk,rst,matrix_A[2928],matrix_B[128],mul_res1[2928]);
multi_7x28 multi_7x28_mod_2929(clk,rst,matrix_A[2929],matrix_B[129],mul_res1[2929]);
multi_7x28 multi_7x28_mod_2930(clk,rst,matrix_A[2930],matrix_B[130],mul_res1[2930]);
multi_7x28 multi_7x28_mod_2931(clk,rst,matrix_A[2931],matrix_B[131],mul_res1[2931]);
multi_7x28 multi_7x28_mod_2932(clk,rst,matrix_A[2932],matrix_B[132],mul_res1[2932]);
multi_7x28 multi_7x28_mod_2933(clk,rst,matrix_A[2933],matrix_B[133],mul_res1[2933]);
multi_7x28 multi_7x28_mod_2934(clk,rst,matrix_A[2934],matrix_B[134],mul_res1[2934]);
multi_7x28 multi_7x28_mod_2935(clk,rst,matrix_A[2935],matrix_B[135],mul_res1[2935]);
multi_7x28 multi_7x28_mod_2936(clk,rst,matrix_A[2936],matrix_B[136],mul_res1[2936]);
multi_7x28 multi_7x28_mod_2937(clk,rst,matrix_A[2937],matrix_B[137],mul_res1[2937]);
multi_7x28 multi_7x28_mod_2938(clk,rst,matrix_A[2938],matrix_B[138],mul_res1[2938]);
multi_7x28 multi_7x28_mod_2939(clk,rst,matrix_A[2939],matrix_B[139],mul_res1[2939]);
multi_7x28 multi_7x28_mod_2940(clk,rst,matrix_A[2940],matrix_B[140],mul_res1[2940]);
multi_7x28 multi_7x28_mod_2941(clk,rst,matrix_A[2941],matrix_B[141],mul_res1[2941]);
multi_7x28 multi_7x28_mod_2942(clk,rst,matrix_A[2942],matrix_B[142],mul_res1[2942]);
multi_7x28 multi_7x28_mod_2943(clk,rst,matrix_A[2943],matrix_B[143],mul_res1[2943]);
multi_7x28 multi_7x28_mod_2944(clk,rst,matrix_A[2944],matrix_B[144],mul_res1[2944]);
multi_7x28 multi_7x28_mod_2945(clk,rst,matrix_A[2945],matrix_B[145],mul_res1[2945]);
multi_7x28 multi_7x28_mod_2946(clk,rst,matrix_A[2946],matrix_B[146],mul_res1[2946]);
multi_7x28 multi_7x28_mod_2947(clk,rst,matrix_A[2947],matrix_B[147],mul_res1[2947]);
multi_7x28 multi_7x28_mod_2948(clk,rst,matrix_A[2948],matrix_B[148],mul_res1[2948]);
multi_7x28 multi_7x28_mod_2949(clk,rst,matrix_A[2949],matrix_B[149],mul_res1[2949]);
multi_7x28 multi_7x28_mod_2950(clk,rst,matrix_A[2950],matrix_B[150],mul_res1[2950]);
multi_7x28 multi_7x28_mod_2951(clk,rst,matrix_A[2951],matrix_B[151],mul_res1[2951]);
multi_7x28 multi_7x28_mod_2952(clk,rst,matrix_A[2952],matrix_B[152],mul_res1[2952]);
multi_7x28 multi_7x28_mod_2953(clk,rst,matrix_A[2953],matrix_B[153],mul_res1[2953]);
multi_7x28 multi_7x28_mod_2954(clk,rst,matrix_A[2954],matrix_B[154],mul_res1[2954]);
multi_7x28 multi_7x28_mod_2955(clk,rst,matrix_A[2955],matrix_B[155],mul_res1[2955]);
multi_7x28 multi_7x28_mod_2956(clk,rst,matrix_A[2956],matrix_B[156],mul_res1[2956]);
multi_7x28 multi_7x28_mod_2957(clk,rst,matrix_A[2957],matrix_B[157],mul_res1[2957]);
multi_7x28 multi_7x28_mod_2958(clk,rst,matrix_A[2958],matrix_B[158],mul_res1[2958]);
multi_7x28 multi_7x28_mod_2959(clk,rst,matrix_A[2959],matrix_B[159],mul_res1[2959]);
multi_7x28 multi_7x28_mod_2960(clk,rst,matrix_A[2960],matrix_B[160],mul_res1[2960]);
multi_7x28 multi_7x28_mod_2961(clk,rst,matrix_A[2961],matrix_B[161],mul_res1[2961]);
multi_7x28 multi_7x28_mod_2962(clk,rst,matrix_A[2962],matrix_B[162],mul_res1[2962]);
multi_7x28 multi_7x28_mod_2963(clk,rst,matrix_A[2963],matrix_B[163],mul_res1[2963]);
multi_7x28 multi_7x28_mod_2964(clk,rst,matrix_A[2964],matrix_B[164],mul_res1[2964]);
multi_7x28 multi_7x28_mod_2965(clk,rst,matrix_A[2965],matrix_B[165],mul_res1[2965]);
multi_7x28 multi_7x28_mod_2966(clk,rst,matrix_A[2966],matrix_B[166],mul_res1[2966]);
multi_7x28 multi_7x28_mod_2967(clk,rst,matrix_A[2967],matrix_B[167],mul_res1[2967]);
multi_7x28 multi_7x28_mod_2968(clk,rst,matrix_A[2968],matrix_B[168],mul_res1[2968]);
multi_7x28 multi_7x28_mod_2969(clk,rst,matrix_A[2969],matrix_B[169],mul_res1[2969]);
multi_7x28 multi_7x28_mod_2970(clk,rst,matrix_A[2970],matrix_B[170],mul_res1[2970]);
multi_7x28 multi_7x28_mod_2971(clk,rst,matrix_A[2971],matrix_B[171],mul_res1[2971]);
multi_7x28 multi_7x28_mod_2972(clk,rst,matrix_A[2972],matrix_B[172],mul_res1[2972]);
multi_7x28 multi_7x28_mod_2973(clk,rst,matrix_A[2973],matrix_B[173],mul_res1[2973]);
multi_7x28 multi_7x28_mod_2974(clk,rst,matrix_A[2974],matrix_B[174],mul_res1[2974]);
multi_7x28 multi_7x28_mod_2975(clk,rst,matrix_A[2975],matrix_B[175],mul_res1[2975]);
multi_7x28 multi_7x28_mod_2976(clk,rst,matrix_A[2976],matrix_B[176],mul_res1[2976]);
multi_7x28 multi_7x28_mod_2977(clk,rst,matrix_A[2977],matrix_B[177],mul_res1[2977]);
multi_7x28 multi_7x28_mod_2978(clk,rst,matrix_A[2978],matrix_B[178],mul_res1[2978]);
multi_7x28 multi_7x28_mod_2979(clk,rst,matrix_A[2979],matrix_B[179],mul_res1[2979]);
multi_7x28 multi_7x28_mod_2980(clk,rst,matrix_A[2980],matrix_B[180],mul_res1[2980]);
multi_7x28 multi_7x28_mod_2981(clk,rst,matrix_A[2981],matrix_B[181],mul_res1[2981]);
multi_7x28 multi_7x28_mod_2982(clk,rst,matrix_A[2982],matrix_B[182],mul_res1[2982]);
multi_7x28 multi_7x28_mod_2983(clk,rst,matrix_A[2983],matrix_B[183],mul_res1[2983]);
multi_7x28 multi_7x28_mod_2984(clk,rst,matrix_A[2984],matrix_B[184],mul_res1[2984]);
multi_7x28 multi_7x28_mod_2985(clk,rst,matrix_A[2985],matrix_B[185],mul_res1[2985]);
multi_7x28 multi_7x28_mod_2986(clk,rst,matrix_A[2986],matrix_B[186],mul_res1[2986]);
multi_7x28 multi_7x28_mod_2987(clk,rst,matrix_A[2987],matrix_B[187],mul_res1[2987]);
multi_7x28 multi_7x28_mod_2988(clk,rst,matrix_A[2988],matrix_B[188],mul_res1[2988]);
multi_7x28 multi_7x28_mod_2989(clk,rst,matrix_A[2989],matrix_B[189],mul_res1[2989]);
multi_7x28 multi_7x28_mod_2990(clk,rst,matrix_A[2990],matrix_B[190],mul_res1[2990]);
multi_7x28 multi_7x28_mod_2991(clk,rst,matrix_A[2991],matrix_B[191],mul_res1[2991]);
multi_7x28 multi_7x28_mod_2992(clk,rst,matrix_A[2992],matrix_B[192],mul_res1[2992]);
multi_7x28 multi_7x28_mod_2993(clk,rst,matrix_A[2993],matrix_B[193],mul_res1[2993]);
multi_7x28 multi_7x28_mod_2994(clk,rst,matrix_A[2994],matrix_B[194],mul_res1[2994]);
multi_7x28 multi_7x28_mod_2995(clk,rst,matrix_A[2995],matrix_B[195],mul_res1[2995]);
multi_7x28 multi_7x28_mod_2996(clk,rst,matrix_A[2996],matrix_B[196],mul_res1[2996]);
multi_7x28 multi_7x28_mod_2997(clk,rst,matrix_A[2997],matrix_B[197],mul_res1[2997]);
multi_7x28 multi_7x28_mod_2998(clk,rst,matrix_A[2998],matrix_B[198],mul_res1[2998]);
multi_7x28 multi_7x28_mod_2999(clk,rst,matrix_A[2999],matrix_B[199],mul_res1[2999]);
multi_7x28 multi_7x28_mod_3000(clk,rst,matrix_A[3000],matrix_B[0],mul_res1[3000]);
multi_7x28 multi_7x28_mod_3001(clk,rst,matrix_A[3001],matrix_B[1],mul_res1[3001]);
multi_7x28 multi_7x28_mod_3002(clk,rst,matrix_A[3002],matrix_B[2],mul_res1[3002]);
multi_7x28 multi_7x28_mod_3003(clk,rst,matrix_A[3003],matrix_B[3],mul_res1[3003]);
multi_7x28 multi_7x28_mod_3004(clk,rst,matrix_A[3004],matrix_B[4],mul_res1[3004]);
multi_7x28 multi_7x28_mod_3005(clk,rst,matrix_A[3005],matrix_B[5],mul_res1[3005]);
multi_7x28 multi_7x28_mod_3006(clk,rst,matrix_A[3006],matrix_B[6],mul_res1[3006]);
multi_7x28 multi_7x28_mod_3007(clk,rst,matrix_A[3007],matrix_B[7],mul_res1[3007]);
multi_7x28 multi_7x28_mod_3008(clk,rst,matrix_A[3008],matrix_B[8],mul_res1[3008]);
multi_7x28 multi_7x28_mod_3009(clk,rst,matrix_A[3009],matrix_B[9],mul_res1[3009]);
multi_7x28 multi_7x28_mod_3010(clk,rst,matrix_A[3010],matrix_B[10],mul_res1[3010]);
multi_7x28 multi_7x28_mod_3011(clk,rst,matrix_A[3011],matrix_B[11],mul_res1[3011]);
multi_7x28 multi_7x28_mod_3012(clk,rst,matrix_A[3012],matrix_B[12],mul_res1[3012]);
multi_7x28 multi_7x28_mod_3013(clk,rst,matrix_A[3013],matrix_B[13],mul_res1[3013]);
multi_7x28 multi_7x28_mod_3014(clk,rst,matrix_A[3014],matrix_B[14],mul_res1[3014]);
multi_7x28 multi_7x28_mod_3015(clk,rst,matrix_A[3015],matrix_B[15],mul_res1[3015]);
multi_7x28 multi_7x28_mod_3016(clk,rst,matrix_A[3016],matrix_B[16],mul_res1[3016]);
multi_7x28 multi_7x28_mod_3017(clk,rst,matrix_A[3017],matrix_B[17],mul_res1[3017]);
multi_7x28 multi_7x28_mod_3018(clk,rst,matrix_A[3018],matrix_B[18],mul_res1[3018]);
multi_7x28 multi_7x28_mod_3019(clk,rst,matrix_A[3019],matrix_B[19],mul_res1[3019]);
multi_7x28 multi_7x28_mod_3020(clk,rst,matrix_A[3020],matrix_B[20],mul_res1[3020]);
multi_7x28 multi_7x28_mod_3021(clk,rst,matrix_A[3021],matrix_B[21],mul_res1[3021]);
multi_7x28 multi_7x28_mod_3022(clk,rst,matrix_A[3022],matrix_B[22],mul_res1[3022]);
multi_7x28 multi_7x28_mod_3023(clk,rst,matrix_A[3023],matrix_B[23],mul_res1[3023]);
multi_7x28 multi_7x28_mod_3024(clk,rst,matrix_A[3024],matrix_B[24],mul_res1[3024]);
multi_7x28 multi_7x28_mod_3025(clk,rst,matrix_A[3025],matrix_B[25],mul_res1[3025]);
multi_7x28 multi_7x28_mod_3026(clk,rst,matrix_A[3026],matrix_B[26],mul_res1[3026]);
multi_7x28 multi_7x28_mod_3027(clk,rst,matrix_A[3027],matrix_B[27],mul_res1[3027]);
multi_7x28 multi_7x28_mod_3028(clk,rst,matrix_A[3028],matrix_B[28],mul_res1[3028]);
multi_7x28 multi_7x28_mod_3029(clk,rst,matrix_A[3029],matrix_B[29],mul_res1[3029]);
multi_7x28 multi_7x28_mod_3030(clk,rst,matrix_A[3030],matrix_B[30],mul_res1[3030]);
multi_7x28 multi_7x28_mod_3031(clk,rst,matrix_A[3031],matrix_B[31],mul_res1[3031]);
multi_7x28 multi_7x28_mod_3032(clk,rst,matrix_A[3032],matrix_B[32],mul_res1[3032]);
multi_7x28 multi_7x28_mod_3033(clk,rst,matrix_A[3033],matrix_B[33],mul_res1[3033]);
multi_7x28 multi_7x28_mod_3034(clk,rst,matrix_A[3034],matrix_B[34],mul_res1[3034]);
multi_7x28 multi_7x28_mod_3035(clk,rst,matrix_A[3035],matrix_B[35],mul_res1[3035]);
multi_7x28 multi_7x28_mod_3036(clk,rst,matrix_A[3036],matrix_B[36],mul_res1[3036]);
multi_7x28 multi_7x28_mod_3037(clk,rst,matrix_A[3037],matrix_B[37],mul_res1[3037]);
multi_7x28 multi_7x28_mod_3038(clk,rst,matrix_A[3038],matrix_B[38],mul_res1[3038]);
multi_7x28 multi_7x28_mod_3039(clk,rst,matrix_A[3039],matrix_B[39],mul_res1[3039]);
multi_7x28 multi_7x28_mod_3040(clk,rst,matrix_A[3040],matrix_B[40],mul_res1[3040]);
multi_7x28 multi_7x28_mod_3041(clk,rst,matrix_A[3041],matrix_B[41],mul_res1[3041]);
multi_7x28 multi_7x28_mod_3042(clk,rst,matrix_A[3042],matrix_B[42],mul_res1[3042]);
multi_7x28 multi_7x28_mod_3043(clk,rst,matrix_A[3043],matrix_B[43],mul_res1[3043]);
multi_7x28 multi_7x28_mod_3044(clk,rst,matrix_A[3044],matrix_B[44],mul_res1[3044]);
multi_7x28 multi_7x28_mod_3045(clk,rst,matrix_A[3045],matrix_B[45],mul_res1[3045]);
multi_7x28 multi_7x28_mod_3046(clk,rst,matrix_A[3046],matrix_B[46],mul_res1[3046]);
multi_7x28 multi_7x28_mod_3047(clk,rst,matrix_A[3047],matrix_B[47],mul_res1[3047]);
multi_7x28 multi_7x28_mod_3048(clk,rst,matrix_A[3048],matrix_B[48],mul_res1[3048]);
multi_7x28 multi_7x28_mod_3049(clk,rst,matrix_A[3049],matrix_B[49],mul_res1[3049]);
multi_7x28 multi_7x28_mod_3050(clk,rst,matrix_A[3050],matrix_B[50],mul_res1[3050]);
multi_7x28 multi_7x28_mod_3051(clk,rst,matrix_A[3051],matrix_B[51],mul_res1[3051]);
multi_7x28 multi_7x28_mod_3052(clk,rst,matrix_A[3052],matrix_B[52],mul_res1[3052]);
multi_7x28 multi_7x28_mod_3053(clk,rst,matrix_A[3053],matrix_B[53],mul_res1[3053]);
multi_7x28 multi_7x28_mod_3054(clk,rst,matrix_A[3054],matrix_B[54],mul_res1[3054]);
multi_7x28 multi_7x28_mod_3055(clk,rst,matrix_A[3055],matrix_B[55],mul_res1[3055]);
multi_7x28 multi_7x28_mod_3056(clk,rst,matrix_A[3056],matrix_B[56],mul_res1[3056]);
multi_7x28 multi_7x28_mod_3057(clk,rst,matrix_A[3057],matrix_B[57],mul_res1[3057]);
multi_7x28 multi_7x28_mod_3058(clk,rst,matrix_A[3058],matrix_B[58],mul_res1[3058]);
multi_7x28 multi_7x28_mod_3059(clk,rst,matrix_A[3059],matrix_B[59],mul_res1[3059]);
multi_7x28 multi_7x28_mod_3060(clk,rst,matrix_A[3060],matrix_B[60],mul_res1[3060]);
multi_7x28 multi_7x28_mod_3061(clk,rst,matrix_A[3061],matrix_B[61],mul_res1[3061]);
multi_7x28 multi_7x28_mod_3062(clk,rst,matrix_A[3062],matrix_B[62],mul_res1[3062]);
multi_7x28 multi_7x28_mod_3063(clk,rst,matrix_A[3063],matrix_B[63],mul_res1[3063]);
multi_7x28 multi_7x28_mod_3064(clk,rst,matrix_A[3064],matrix_B[64],mul_res1[3064]);
multi_7x28 multi_7x28_mod_3065(clk,rst,matrix_A[3065],matrix_B[65],mul_res1[3065]);
multi_7x28 multi_7x28_mod_3066(clk,rst,matrix_A[3066],matrix_B[66],mul_res1[3066]);
multi_7x28 multi_7x28_mod_3067(clk,rst,matrix_A[3067],matrix_B[67],mul_res1[3067]);
multi_7x28 multi_7x28_mod_3068(clk,rst,matrix_A[3068],matrix_B[68],mul_res1[3068]);
multi_7x28 multi_7x28_mod_3069(clk,rst,matrix_A[3069],matrix_B[69],mul_res1[3069]);
multi_7x28 multi_7x28_mod_3070(clk,rst,matrix_A[3070],matrix_B[70],mul_res1[3070]);
multi_7x28 multi_7x28_mod_3071(clk,rst,matrix_A[3071],matrix_B[71],mul_res1[3071]);
multi_7x28 multi_7x28_mod_3072(clk,rst,matrix_A[3072],matrix_B[72],mul_res1[3072]);
multi_7x28 multi_7x28_mod_3073(clk,rst,matrix_A[3073],matrix_B[73],mul_res1[3073]);
multi_7x28 multi_7x28_mod_3074(clk,rst,matrix_A[3074],matrix_B[74],mul_res1[3074]);
multi_7x28 multi_7x28_mod_3075(clk,rst,matrix_A[3075],matrix_B[75],mul_res1[3075]);
multi_7x28 multi_7x28_mod_3076(clk,rst,matrix_A[3076],matrix_B[76],mul_res1[3076]);
multi_7x28 multi_7x28_mod_3077(clk,rst,matrix_A[3077],matrix_B[77],mul_res1[3077]);
multi_7x28 multi_7x28_mod_3078(clk,rst,matrix_A[3078],matrix_B[78],mul_res1[3078]);
multi_7x28 multi_7x28_mod_3079(clk,rst,matrix_A[3079],matrix_B[79],mul_res1[3079]);
multi_7x28 multi_7x28_mod_3080(clk,rst,matrix_A[3080],matrix_B[80],mul_res1[3080]);
multi_7x28 multi_7x28_mod_3081(clk,rst,matrix_A[3081],matrix_B[81],mul_res1[3081]);
multi_7x28 multi_7x28_mod_3082(clk,rst,matrix_A[3082],matrix_B[82],mul_res1[3082]);
multi_7x28 multi_7x28_mod_3083(clk,rst,matrix_A[3083],matrix_B[83],mul_res1[3083]);
multi_7x28 multi_7x28_mod_3084(clk,rst,matrix_A[3084],matrix_B[84],mul_res1[3084]);
multi_7x28 multi_7x28_mod_3085(clk,rst,matrix_A[3085],matrix_B[85],mul_res1[3085]);
multi_7x28 multi_7x28_mod_3086(clk,rst,matrix_A[3086],matrix_B[86],mul_res1[3086]);
multi_7x28 multi_7x28_mod_3087(clk,rst,matrix_A[3087],matrix_B[87],mul_res1[3087]);
multi_7x28 multi_7x28_mod_3088(clk,rst,matrix_A[3088],matrix_B[88],mul_res1[3088]);
multi_7x28 multi_7x28_mod_3089(clk,rst,matrix_A[3089],matrix_B[89],mul_res1[3089]);
multi_7x28 multi_7x28_mod_3090(clk,rst,matrix_A[3090],matrix_B[90],mul_res1[3090]);
multi_7x28 multi_7x28_mod_3091(clk,rst,matrix_A[3091],matrix_B[91],mul_res1[3091]);
multi_7x28 multi_7x28_mod_3092(clk,rst,matrix_A[3092],matrix_B[92],mul_res1[3092]);
multi_7x28 multi_7x28_mod_3093(clk,rst,matrix_A[3093],matrix_B[93],mul_res1[3093]);
multi_7x28 multi_7x28_mod_3094(clk,rst,matrix_A[3094],matrix_B[94],mul_res1[3094]);
multi_7x28 multi_7x28_mod_3095(clk,rst,matrix_A[3095],matrix_B[95],mul_res1[3095]);
multi_7x28 multi_7x28_mod_3096(clk,rst,matrix_A[3096],matrix_B[96],mul_res1[3096]);
multi_7x28 multi_7x28_mod_3097(clk,rst,matrix_A[3097],matrix_B[97],mul_res1[3097]);
multi_7x28 multi_7x28_mod_3098(clk,rst,matrix_A[3098],matrix_B[98],mul_res1[3098]);
multi_7x28 multi_7x28_mod_3099(clk,rst,matrix_A[3099],matrix_B[99],mul_res1[3099]);
multi_7x28 multi_7x28_mod_3100(clk,rst,matrix_A[3100],matrix_B[100],mul_res1[3100]);
multi_7x28 multi_7x28_mod_3101(clk,rst,matrix_A[3101],matrix_B[101],mul_res1[3101]);
multi_7x28 multi_7x28_mod_3102(clk,rst,matrix_A[3102],matrix_B[102],mul_res1[3102]);
multi_7x28 multi_7x28_mod_3103(clk,rst,matrix_A[3103],matrix_B[103],mul_res1[3103]);
multi_7x28 multi_7x28_mod_3104(clk,rst,matrix_A[3104],matrix_B[104],mul_res1[3104]);
multi_7x28 multi_7x28_mod_3105(clk,rst,matrix_A[3105],matrix_B[105],mul_res1[3105]);
multi_7x28 multi_7x28_mod_3106(clk,rst,matrix_A[3106],matrix_B[106],mul_res1[3106]);
multi_7x28 multi_7x28_mod_3107(clk,rst,matrix_A[3107],matrix_B[107],mul_res1[3107]);
multi_7x28 multi_7x28_mod_3108(clk,rst,matrix_A[3108],matrix_B[108],mul_res1[3108]);
multi_7x28 multi_7x28_mod_3109(clk,rst,matrix_A[3109],matrix_B[109],mul_res1[3109]);
multi_7x28 multi_7x28_mod_3110(clk,rst,matrix_A[3110],matrix_B[110],mul_res1[3110]);
multi_7x28 multi_7x28_mod_3111(clk,rst,matrix_A[3111],matrix_B[111],mul_res1[3111]);
multi_7x28 multi_7x28_mod_3112(clk,rst,matrix_A[3112],matrix_B[112],mul_res1[3112]);
multi_7x28 multi_7x28_mod_3113(clk,rst,matrix_A[3113],matrix_B[113],mul_res1[3113]);
multi_7x28 multi_7x28_mod_3114(clk,rst,matrix_A[3114],matrix_B[114],mul_res1[3114]);
multi_7x28 multi_7x28_mod_3115(clk,rst,matrix_A[3115],matrix_B[115],mul_res1[3115]);
multi_7x28 multi_7x28_mod_3116(clk,rst,matrix_A[3116],matrix_B[116],mul_res1[3116]);
multi_7x28 multi_7x28_mod_3117(clk,rst,matrix_A[3117],matrix_B[117],mul_res1[3117]);
multi_7x28 multi_7x28_mod_3118(clk,rst,matrix_A[3118],matrix_B[118],mul_res1[3118]);
multi_7x28 multi_7x28_mod_3119(clk,rst,matrix_A[3119],matrix_B[119],mul_res1[3119]);
multi_7x28 multi_7x28_mod_3120(clk,rst,matrix_A[3120],matrix_B[120],mul_res1[3120]);
multi_7x28 multi_7x28_mod_3121(clk,rst,matrix_A[3121],matrix_B[121],mul_res1[3121]);
multi_7x28 multi_7x28_mod_3122(clk,rst,matrix_A[3122],matrix_B[122],mul_res1[3122]);
multi_7x28 multi_7x28_mod_3123(clk,rst,matrix_A[3123],matrix_B[123],mul_res1[3123]);
multi_7x28 multi_7x28_mod_3124(clk,rst,matrix_A[3124],matrix_B[124],mul_res1[3124]);
multi_7x28 multi_7x28_mod_3125(clk,rst,matrix_A[3125],matrix_B[125],mul_res1[3125]);
multi_7x28 multi_7x28_mod_3126(clk,rst,matrix_A[3126],matrix_B[126],mul_res1[3126]);
multi_7x28 multi_7x28_mod_3127(clk,rst,matrix_A[3127],matrix_B[127],mul_res1[3127]);
multi_7x28 multi_7x28_mod_3128(clk,rst,matrix_A[3128],matrix_B[128],mul_res1[3128]);
multi_7x28 multi_7x28_mod_3129(clk,rst,matrix_A[3129],matrix_B[129],mul_res1[3129]);
multi_7x28 multi_7x28_mod_3130(clk,rst,matrix_A[3130],matrix_B[130],mul_res1[3130]);
multi_7x28 multi_7x28_mod_3131(clk,rst,matrix_A[3131],matrix_B[131],mul_res1[3131]);
multi_7x28 multi_7x28_mod_3132(clk,rst,matrix_A[3132],matrix_B[132],mul_res1[3132]);
multi_7x28 multi_7x28_mod_3133(clk,rst,matrix_A[3133],matrix_B[133],mul_res1[3133]);
multi_7x28 multi_7x28_mod_3134(clk,rst,matrix_A[3134],matrix_B[134],mul_res1[3134]);
multi_7x28 multi_7x28_mod_3135(clk,rst,matrix_A[3135],matrix_B[135],mul_res1[3135]);
multi_7x28 multi_7x28_mod_3136(clk,rst,matrix_A[3136],matrix_B[136],mul_res1[3136]);
multi_7x28 multi_7x28_mod_3137(clk,rst,matrix_A[3137],matrix_B[137],mul_res1[3137]);
multi_7x28 multi_7x28_mod_3138(clk,rst,matrix_A[3138],matrix_B[138],mul_res1[3138]);
multi_7x28 multi_7x28_mod_3139(clk,rst,matrix_A[3139],matrix_B[139],mul_res1[3139]);
multi_7x28 multi_7x28_mod_3140(clk,rst,matrix_A[3140],matrix_B[140],mul_res1[3140]);
multi_7x28 multi_7x28_mod_3141(clk,rst,matrix_A[3141],matrix_B[141],mul_res1[3141]);
multi_7x28 multi_7x28_mod_3142(clk,rst,matrix_A[3142],matrix_B[142],mul_res1[3142]);
multi_7x28 multi_7x28_mod_3143(clk,rst,matrix_A[3143],matrix_B[143],mul_res1[3143]);
multi_7x28 multi_7x28_mod_3144(clk,rst,matrix_A[3144],matrix_B[144],mul_res1[3144]);
multi_7x28 multi_7x28_mod_3145(clk,rst,matrix_A[3145],matrix_B[145],mul_res1[3145]);
multi_7x28 multi_7x28_mod_3146(clk,rst,matrix_A[3146],matrix_B[146],mul_res1[3146]);
multi_7x28 multi_7x28_mod_3147(clk,rst,matrix_A[3147],matrix_B[147],mul_res1[3147]);
multi_7x28 multi_7x28_mod_3148(clk,rst,matrix_A[3148],matrix_B[148],mul_res1[3148]);
multi_7x28 multi_7x28_mod_3149(clk,rst,matrix_A[3149],matrix_B[149],mul_res1[3149]);
multi_7x28 multi_7x28_mod_3150(clk,rst,matrix_A[3150],matrix_B[150],mul_res1[3150]);
multi_7x28 multi_7x28_mod_3151(clk,rst,matrix_A[3151],matrix_B[151],mul_res1[3151]);
multi_7x28 multi_7x28_mod_3152(clk,rst,matrix_A[3152],matrix_B[152],mul_res1[3152]);
multi_7x28 multi_7x28_mod_3153(clk,rst,matrix_A[3153],matrix_B[153],mul_res1[3153]);
multi_7x28 multi_7x28_mod_3154(clk,rst,matrix_A[3154],matrix_B[154],mul_res1[3154]);
multi_7x28 multi_7x28_mod_3155(clk,rst,matrix_A[3155],matrix_B[155],mul_res1[3155]);
multi_7x28 multi_7x28_mod_3156(clk,rst,matrix_A[3156],matrix_B[156],mul_res1[3156]);
multi_7x28 multi_7x28_mod_3157(clk,rst,matrix_A[3157],matrix_B[157],mul_res1[3157]);
multi_7x28 multi_7x28_mod_3158(clk,rst,matrix_A[3158],matrix_B[158],mul_res1[3158]);
multi_7x28 multi_7x28_mod_3159(clk,rst,matrix_A[3159],matrix_B[159],mul_res1[3159]);
multi_7x28 multi_7x28_mod_3160(clk,rst,matrix_A[3160],matrix_B[160],mul_res1[3160]);
multi_7x28 multi_7x28_mod_3161(clk,rst,matrix_A[3161],matrix_B[161],mul_res1[3161]);
multi_7x28 multi_7x28_mod_3162(clk,rst,matrix_A[3162],matrix_B[162],mul_res1[3162]);
multi_7x28 multi_7x28_mod_3163(clk,rst,matrix_A[3163],matrix_B[163],mul_res1[3163]);
multi_7x28 multi_7x28_mod_3164(clk,rst,matrix_A[3164],matrix_B[164],mul_res1[3164]);
multi_7x28 multi_7x28_mod_3165(clk,rst,matrix_A[3165],matrix_B[165],mul_res1[3165]);
multi_7x28 multi_7x28_mod_3166(clk,rst,matrix_A[3166],matrix_B[166],mul_res1[3166]);
multi_7x28 multi_7x28_mod_3167(clk,rst,matrix_A[3167],matrix_B[167],mul_res1[3167]);
multi_7x28 multi_7x28_mod_3168(clk,rst,matrix_A[3168],matrix_B[168],mul_res1[3168]);
multi_7x28 multi_7x28_mod_3169(clk,rst,matrix_A[3169],matrix_B[169],mul_res1[3169]);
multi_7x28 multi_7x28_mod_3170(clk,rst,matrix_A[3170],matrix_B[170],mul_res1[3170]);
multi_7x28 multi_7x28_mod_3171(clk,rst,matrix_A[3171],matrix_B[171],mul_res1[3171]);
multi_7x28 multi_7x28_mod_3172(clk,rst,matrix_A[3172],matrix_B[172],mul_res1[3172]);
multi_7x28 multi_7x28_mod_3173(clk,rst,matrix_A[3173],matrix_B[173],mul_res1[3173]);
multi_7x28 multi_7x28_mod_3174(clk,rst,matrix_A[3174],matrix_B[174],mul_res1[3174]);
multi_7x28 multi_7x28_mod_3175(clk,rst,matrix_A[3175],matrix_B[175],mul_res1[3175]);
multi_7x28 multi_7x28_mod_3176(clk,rst,matrix_A[3176],matrix_B[176],mul_res1[3176]);
multi_7x28 multi_7x28_mod_3177(clk,rst,matrix_A[3177],matrix_B[177],mul_res1[3177]);
multi_7x28 multi_7x28_mod_3178(clk,rst,matrix_A[3178],matrix_B[178],mul_res1[3178]);
multi_7x28 multi_7x28_mod_3179(clk,rst,matrix_A[3179],matrix_B[179],mul_res1[3179]);
multi_7x28 multi_7x28_mod_3180(clk,rst,matrix_A[3180],matrix_B[180],mul_res1[3180]);
multi_7x28 multi_7x28_mod_3181(clk,rst,matrix_A[3181],matrix_B[181],mul_res1[3181]);
multi_7x28 multi_7x28_mod_3182(clk,rst,matrix_A[3182],matrix_B[182],mul_res1[3182]);
multi_7x28 multi_7x28_mod_3183(clk,rst,matrix_A[3183],matrix_B[183],mul_res1[3183]);
multi_7x28 multi_7x28_mod_3184(clk,rst,matrix_A[3184],matrix_B[184],mul_res1[3184]);
multi_7x28 multi_7x28_mod_3185(clk,rst,matrix_A[3185],matrix_B[185],mul_res1[3185]);
multi_7x28 multi_7x28_mod_3186(clk,rst,matrix_A[3186],matrix_B[186],mul_res1[3186]);
multi_7x28 multi_7x28_mod_3187(clk,rst,matrix_A[3187],matrix_B[187],mul_res1[3187]);
multi_7x28 multi_7x28_mod_3188(clk,rst,matrix_A[3188],matrix_B[188],mul_res1[3188]);
multi_7x28 multi_7x28_mod_3189(clk,rst,matrix_A[3189],matrix_B[189],mul_res1[3189]);
multi_7x28 multi_7x28_mod_3190(clk,rst,matrix_A[3190],matrix_B[190],mul_res1[3190]);
multi_7x28 multi_7x28_mod_3191(clk,rst,matrix_A[3191],matrix_B[191],mul_res1[3191]);
multi_7x28 multi_7x28_mod_3192(clk,rst,matrix_A[3192],matrix_B[192],mul_res1[3192]);
multi_7x28 multi_7x28_mod_3193(clk,rst,matrix_A[3193],matrix_B[193],mul_res1[3193]);
multi_7x28 multi_7x28_mod_3194(clk,rst,matrix_A[3194],matrix_B[194],mul_res1[3194]);
multi_7x28 multi_7x28_mod_3195(clk,rst,matrix_A[3195],matrix_B[195],mul_res1[3195]);
multi_7x28 multi_7x28_mod_3196(clk,rst,matrix_A[3196],matrix_B[196],mul_res1[3196]);
multi_7x28 multi_7x28_mod_3197(clk,rst,matrix_A[3197],matrix_B[197],mul_res1[3197]);
multi_7x28 multi_7x28_mod_3198(clk,rst,matrix_A[3198],matrix_B[198],mul_res1[3198]);
multi_7x28 multi_7x28_mod_3199(clk,rst,matrix_A[3199],matrix_B[199],mul_res1[3199]);
multi_7x28 multi_7x28_mod_3200(clk,rst,matrix_A[3200],matrix_B[0],mul_res1[3200]);
multi_7x28 multi_7x28_mod_3201(clk,rst,matrix_A[3201],matrix_B[1],mul_res1[3201]);
multi_7x28 multi_7x28_mod_3202(clk,rst,matrix_A[3202],matrix_B[2],mul_res1[3202]);
multi_7x28 multi_7x28_mod_3203(clk,rst,matrix_A[3203],matrix_B[3],mul_res1[3203]);
multi_7x28 multi_7x28_mod_3204(clk,rst,matrix_A[3204],matrix_B[4],mul_res1[3204]);
multi_7x28 multi_7x28_mod_3205(clk,rst,matrix_A[3205],matrix_B[5],mul_res1[3205]);
multi_7x28 multi_7x28_mod_3206(clk,rst,matrix_A[3206],matrix_B[6],mul_res1[3206]);
multi_7x28 multi_7x28_mod_3207(clk,rst,matrix_A[3207],matrix_B[7],mul_res1[3207]);
multi_7x28 multi_7x28_mod_3208(clk,rst,matrix_A[3208],matrix_B[8],mul_res1[3208]);
multi_7x28 multi_7x28_mod_3209(clk,rst,matrix_A[3209],matrix_B[9],mul_res1[3209]);
multi_7x28 multi_7x28_mod_3210(clk,rst,matrix_A[3210],matrix_B[10],mul_res1[3210]);
multi_7x28 multi_7x28_mod_3211(clk,rst,matrix_A[3211],matrix_B[11],mul_res1[3211]);
multi_7x28 multi_7x28_mod_3212(clk,rst,matrix_A[3212],matrix_B[12],mul_res1[3212]);
multi_7x28 multi_7x28_mod_3213(clk,rst,matrix_A[3213],matrix_B[13],mul_res1[3213]);
multi_7x28 multi_7x28_mod_3214(clk,rst,matrix_A[3214],matrix_B[14],mul_res1[3214]);
multi_7x28 multi_7x28_mod_3215(clk,rst,matrix_A[3215],matrix_B[15],mul_res1[3215]);
multi_7x28 multi_7x28_mod_3216(clk,rst,matrix_A[3216],matrix_B[16],mul_res1[3216]);
multi_7x28 multi_7x28_mod_3217(clk,rst,matrix_A[3217],matrix_B[17],mul_res1[3217]);
multi_7x28 multi_7x28_mod_3218(clk,rst,matrix_A[3218],matrix_B[18],mul_res1[3218]);
multi_7x28 multi_7x28_mod_3219(clk,rst,matrix_A[3219],matrix_B[19],mul_res1[3219]);
multi_7x28 multi_7x28_mod_3220(clk,rst,matrix_A[3220],matrix_B[20],mul_res1[3220]);
multi_7x28 multi_7x28_mod_3221(clk,rst,matrix_A[3221],matrix_B[21],mul_res1[3221]);
multi_7x28 multi_7x28_mod_3222(clk,rst,matrix_A[3222],matrix_B[22],mul_res1[3222]);
multi_7x28 multi_7x28_mod_3223(clk,rst,matrix_A[3223],matrix_B[23],mul_res1[3223]);
multi_7x28 multi_7x28_mod_3224(clk,rst,matrix_A[3224],matrix_B[24],mul_res1[3224]);
multi_7x28 multi_7x28_mod_3225(clk,rst,matrix_A[3225],matrix_B[25],mul_res1[3225]);
multi_7x28 multi_7x28_mod_3226(clk,rst,matrix_A[3226],matrix_B[26],mul_res1[3226]);
multi_7x28 multi_7x28_mod_3227(clk,rst,matrix_A[3227],matrix_B[27],mul_res1[3227]);
multi_7x28 multi_7x28_mod_3228(clk,rst,matrix_A[3228],matrix_B[28],mul_res1[3228]);
multi_7x28 multi_7x28_mod_3229(clk,rst,matrix_A[3229],matrix_B[29],mul_res1[3229]);
multi_7x28 multi_7x28_mod_3230(clk,rst,matrix_A[3230],matrix_B[30],mul_res1[3230]);
multi_7x28 multi_7x28_mod_3231(clk,rst,matrix_A[3231],matrix_B[31],mul_res1[3231]);
multi_7x28 multi_7x28_mod_3232(clk,rst,matrix_A[3232],matrix_B[32],mul_res1[3232]);
multi_7x28 multi_7x28_mod_3233(clk,rst,matrix_A[3233],matrix_B[33],mul_res1[3233]);
multi_7x28 multi_7x28_mod_3234(clk,rst,matrix_A[3234],matrix_B[34],mul_res1[3234]);
multi_7x28 multi_7x28_mod_3235(clk,rst,matrix_A[3235],matrix_B[35],mul_res1[3235]);
multi_7x28 multi_7x28_mod_3236(clk,rst,matrix_A[3236],matrix_B[36],mul_res1[3236]);
multi_7x28 multi_7x28_mod_3237(clk,rst,matrix_A[3237],matrix_B[37],mul_res1[3237]);
multi_7x28 multi_7x28_mod_3238(clk,rst,matrix_A[3238],matrix_B[38],mul_res1[3238]);
multi_7x28 multi_7x28_mod_3239(clk,rst,matrix_A[3239],matrix_B[39],mul_res1[3239]);
multi_7x28 multi_7x28_mod_3240(clk,rst,matrix_A[3240],matrix_B[40],mul_res1[3240]);
multi_7x28 multi_7x28_mod_3241(clk,rst,matrix_A[3241],matrix_B[41],mul_res1[3241]);
multi_7x28 multi_7x28_mod_3242(clk,rst,matrix_A[3242],matrix_B[42],mul_res1[3242]);
multi_7x28 multi_7x28_mod_3243(clk,rst,matrix_A[3243],matrix_B[43],mul_res1[3243]);
multi_7x28 multi_7x28_mod_3244(clk,rst,matrix_A[3244],matrix_B[44],mul_res1[3244]);
multi_7x28 multi_7x28_mod_3245(clk,rst,matrix_A[3245],matrix_B[45],mul_res1[3245]);
multi_7x28 multi_7x28_mod_3246(clk,rst,matrix_A[3246],matrix_B[46],mul_res1[3246]);
multi_7x28 multi_7x28_mod_3247(clk,rst,matrix_A[3247],matrix_B[47],mul_res1[3247]);
multi_7x28 multi_7x28_mod_3248(clk,rst,matrix_A[3248],matrix_B[48],mul_res1[3248]);
multi_7x28 multi_7x28_mod_3249(clk,rst,matrix_A[3249],matrix_B[49],mul_res1[3249]);
multi_7x28 multi_7x28_mod_3250(clk,rst,matrix_A[3250],matrix_B[50],mul_res1[3250]);
multi_7x28 multi_7x28_mod_3251(clk,rst,matrix_A[3251],matrix_B[51],mul_res1[3251]);
multi_7x28 multi_7x28_mod_3252(clk,rst,matrix_A[3252],matrix_B[52],mul_res1[3252]);
multi_7x28 multi_7x28_mod_3253(clk,rst,matrix_A[3253],matrix_B[53],mul_res1[3253]);
multi_7x28 multi_7x28_mod_3254(clk,rst,matrix_A[3254],matrix_B[54],mul_res1[3254]);
multi_7x28 multi_7x28_mod_3255(clk,rst,matrix_A[3255],matrix_B[55],mul_res1[3255]);
multi_7x28 multi_7x28_mod_3256(clk,rst,matrix_A[3256],matrix_B[56],mul_res1[3256]);
multi_7x28 multi_7x28_mod_3257(clk,rst,matrix_A[3257],matrix_B[57],mul_res1[3257]);
multi_7x28 multi_7x28_mod_3258(clk,rst,matrix_A[3258],matrix_B[58],mul_res1[3258]);
multi_7x28 multi_7x28_mod_3259(clk,rst,matrix_A[3259],matrix_B[59],mul_res1[3259]);
multi_7x28 multi_7x28_mod_3260(clk,rst,matrix_A[3260],matrix_B[60],mul_res1[3260]);
multi_7x28 multi_7x28_mod_3261(clk,rst,matrix_A[3261],matrix_B[61],mul_res1[3261]);
multi_7x28 multi_7x28_mod_3262(clk,rst,matrix_A[3262],matrix_B[62],mul_res1[3262]);
multi_7x28 multi_7x28_mod_3263(clk,rst,matrix_A[3263],matrix_B[63],mul_res1[3263]);
multi_7x28 multi_7x28_mod_3264(clk,rst,matrix_A[3264],matrix_B[64],mul_res1[3264]);
multi_7x28 multi_7x28_mod_3265(clk,rst,matrix_A[3265],matrix_B[65],mul_res1[3265]);
multi_7x28 multi_7x28_mod_3266(clk,rst,matrix_A[3266],matrix_B[66],mul_res1[3266]);
multi_7x28 multi_7x28_mod_3267(clk,rst,matrix_A[3267],matrix_B[67],mul_res1[3267]);
multi_7x28 multi_7x28_mod_3268(clk,rst,matrix_A[3268],matrix_B[68],mul_res1[3268]);
multi_7x28 multi_7x28_mod_3269(clk,rst,matrix_A[3269],matrix_B[69],mul_res1[3269]);
multi_7x28 multi_7x28_mod_3270(clk,rst,matrix_A[3270],matrix_B[70],mul_res1[3270]);
multi_7x28 multi_7x28_mod_3271(clk,rst,matrix_A[3271],matrix_B[71],mul_res1[3271]);
multi_7x28 multi_7x28_mod_3272(clk,rst,matrix_A[3272],matrix_B[72],mul_res1[3272]);
multi_7x28 multi_7x28_mod_3273(clk,rst,matrix_A[3273],matrix_B[73],mul_res1[3273]);
multi_7x28 multi_7x28_mod_3274(clk,rst,matrix_A[3274],matrix_B[74],mul_res1[3274]);
multi_7x28 multi_7x28_mod_3275(clk,rst,matrix_A[3275],matrix_B[75],mul_res1[3275]);
multi_7x28 multi_7x28_mod_3276(clk,rst,matrix_A[3276],matrix_B[76],mul_res1[3276]);
multi_7x28 multi_7x28_mod_3277(clk,rst,matrix_A[3277],matrix_B[77],mul_res1[3277]);
multi_7x28 multi_7x28_mod_3278(clk,rst,matrix_A[3278],matrix_B[78],mul_res1[3278]);
multi_7x28 multi_7x28_mod_3279(clk,rst,matrix_A[3279],matrix_B[79],mul_res1[3279]);
multi_7x28 multi_7x28_mod_3280(clk,rst,matrix_A[3280],matrix_B[80],mul_res1[3280]);
multi_7x28 multi_7x28_mod_3281(clk,rst,matrix_A[3281],matrix_B[81],mul_res1[3281]);
multi_7x28 multi_7x28_mod_3282(clk,rst,matrix_A[3282],matrix_B[82],mul_res1[3282]);
multi_7x28 multi_7x28_mod_3283(clk,rst,matrix_A[3283],matrix_B[83],mul_res1[3283]);
multi_7x28 multi_7x28_mod_3284(clk,rst,matrix_A[3284],matrix_B[84],mul_res1[3284]);
multi_7x28 multi_7x28_mod_3285(clk,rst,matrix_A[3285],matrix_B[85],mul_res1[3285]);
multi_7x28 multi_7x28_mod_3286(clk,rst,matrix_A[3286],matrix_B[86],mul_res1[3286]);
multi_7x28 multi_7x28_mod_3287(clk,rst,matrix_A[3287],matrix_B[87],mul_res1[3287]);
multi_7x28 multi_7x28_mod_3288(clk,rst,matrix_A[3288],matrix_B[88],mul_res1[3288]);
multi_7x28 multi_7x28_mod_3289(clk,rst,matrix_A[3289],matrix_B[89],mul_res1[3289]);
multi_7x28 multi_7x28_mod_3290(clk,rst,matrix_A[3290],matrix_B[90],mul_res1[3290]);
multi_7x28 multi_7x28_mod_3291(clk,rst,matrix_A[3291],matrix_B[91],mul_res1[3291]);
multi_7x28 multi_7x28_mod_3292(clk,rst,matrix_A[3292],matrix_B[92],mul_res1[3292]);
multi_7x28 multi_7x28_mod_3293(clk,rst,matrix_A[3293],matrix_B[93],mul_res1[3293]);
multi_7x28 multi_7x28_mod_3294(clk,rst,matrix_A[3294],matrix_B[94],mul_res1[3294]);
multi_7x28 multi_7x28_mod_3295(clk,rst,matrix_A[3295],matrix_B[95],mul_res1[3295]);
multi_7x28 multi_7x28_mod_3296(clk,rst,matrix_A[3296],matrix_B[96],mul_res1[3296]);
multi_7x28 multi_7x28_mod_3297(clk,rst,matrix_A[3297],matrix_B[97],mul_res1[3297]);
multi_7x28 multi_7x28_mod_3298(clk,rst,matrix_A[3298],matrix_B[98],mul_res1[3298]);
multi_7x28 multi_7x28_mod_3299(clk,rst,matrix_A[3299],matrix_B[99],mul_res1[3299]);
multi_7x28 multi_7x28_mod_3300(clk,rst,matrix_A[3300],matrix_B[100],mul_res1[3300]);
multi_7x28 multi_7x28_mod_3301(clk,rst,matrix_A[3301],matrix_B[101],mul_res1[3301]);
multi_7x28 multi_7x28_mod_3302(clk,rst,matrix_A[3302],matrix_B[102],mul_res1[3302]);
multi_7x28 multi_7x28_mod_3303(clk,rst,matrix_A[3303],matrix_B[103],mul_res1[3303]);
multi_7x28 multi_7x28_mod_3304(clk,rst,matrix_A[3304],matrix_B[104],mul_res1[3304]);
multi_7x28 multi_7x28_mod_3305(clk,rst,matrix_A[3305],matrix_B[105],mul_res1[3305]);
multi_7x28 multi_7x28_mod_3306(clk,rst,matrix_A[3306],matrix_B[106],mul_res1[3306]);
multi_7x28 multi_7x28_mod_3307(clk,rst,matrix_A[3307],matrix_B[107],mul_res1[3307]);
multi_7x28 multi_7x28_mod_3308(clk,rst,matrix_A[3308],matrix_B[108],mul_res1[3308]);
multi_7x28 multi_7x28_mod_3309(clk,rst,matrix_A[3309],matrix_B[109],mul_res1[3309]);
multi_7x28 multi_7x28_mod_3310(clk,rst,matrix_A[3310],matrix_B[110],mul_res1[3310]);
multi_7x28 multi_7x28_mod_3311(clk,rst,matrix_A[3311],matrix_B[111],mul_res1[3311]);
multi_7x28 multi_7x28_mod_3312(clk,rst,matrix_A[3312],matrix_B[112],mul_res1[3312]);
multi_7x28 multi_7x28_mod_3313(clk,rst,matrix_A[3313],matrix_B[113],mul_res1[3313]);
multi_7x28 multi_7x28_mod_3314(clk,rst,matrix_A[3314],matrix_B[114],mul_res1[3314]);
multi_7x28 multi_7x28_mod_3315(clk,rst,matrix_A[3315],matrix_B[115],mul_res1[3315]);
multi_7x28 multi_7x28_mod_3316(clk,rst,matrix_A[3316],matrix_B[116],mul_res1[3316]);
multi_7x28 multi_7x28_mod_3317(clk,rst,matrix_A[3317],matrix_B[117],mul_res1[3317]);
multi_7x28 multi_7x28_mod_3318(clk,rst,matrix_A[3318],matrix_B[118],mul_res1[3318]);
multi_7x28 multi_7x28_mod_3319(clk,rst,matrix_A[3319],matrix_B[119],mul_res1[3319]);
multi_7x28 multi_7x28_mod_3320(clk,rst,matrix_A[3320],matrix_B[120],mul_res1[3320]);
multi_7x28 multi_7x28_mod_3321(clk,rst,matrix_A[3321],matrix_B[121],mul_res1[3321]);
multi_7x28 multi_7x28_mod_3322(clk,rst,matrix_A[3322],matrix_B[122],mul_res1[3322]);
multi_7x28 multi_7x28_mod_3323(clk,rst,matrix_A[3323],matrix_B[123],mul_res1[3323]);
multi_7x28 multi_7x28_mod_3324(clk,rst,matrix_A[3324],matrix_B[124],mul_res1[3324]);
multi_7x28 multi_7x28_mod_3325(clk,rst,matrix_A[3325],matrix_B[125],mul_res1[3325]);
multi_7x28 multi_7x28_mod_3326(clk,rst,matrix_A[3326],matrix_B[126],mul_res1[3326]);
multi_7x28 multi_7x28_mod_3327(clk,rst,matrix_A[3327],matrix_B[127],mul_res1[3327]);
multi_7x28 multi_7x28_mod_3328(clk,rst,matrix_A[3328],matrix_B[128],mul_res1[3328]);
multi_7x28 multi_7x28_mod_3329(clk,rst,matrix_A[3329],matrix_B[129],mul_res1[3329]);
multi_7x28 multi_7x28_mod_3330(clk,rst,matrix_A[3330],matrix_B[130],mul_res1[3330]);
multi_7x28 multi_7x28_mod_3331(clk,rst,matrix_A[3331],matrix_B[131],mul_res1[3331]);
multi_7x28 multi_7x28_mod_3332(clk,rst,matrix_A[3332],matrix_B[132],mul_res1[3332]);
multi_7x28 multi_7x28_mod_3333(clk,rst,matrix_A[3333],matrix_B[133],mul_res1[3333]);
multi_7x28 multi_7x28_mod_3334(clk,rst,matrix_A[3334],matrix_B[134],mul_res1[3334]);
multi_7x28 multi_7x28_mod_3335(clk,rst,matrix_A[3335],matrix_B[135],mul_res1[3335]);
multi_7x28 multi_7x28_mod_3336(clk,rst,matrix_A[3336],matrix_B[136],mul_res1[3336]);
multi_7x28 multi_7x28_mod_3337(clk,rst,matrix_A[3337],matrix_B[137],mul_res1[3337]);
multi_7x28 multi_7x28_mod_3338(clk,rst,matrix_A[3338],matrix_B[138],mul_res1[3338]);
multi_7x28 multi_7x28_mod_3339(clk,rst,matrix_A[3339],matrix_B[139],mul_res1[3339]);
multi_7x28 multi_7x28_mod_3340(clk,rst,matrix_A[3340],matrix_B[140],mul_res1[3340]);
multi_7x28 multi_7x28_mod_3341(clk,rst,matrix_A[3341],matrix_B[141],mul_res1[3341]);
multi_7x28 multi_7x28_mod_3342(clk,rst,matrix_A[3342],matrix_B[142],mul_res1[3342]);
multi_7x28 multi_7x28_mod_3343(clk,rst,matrix_A[3343],matrix_B[143],mul_res1[3343]);
multi_7x28 multi_7x28_mod_3344(clk,rst,matrix_A[3344],matrix_B[144],mul_res1[3344]);
multi_7x28 multi_7x28_mod_3345(clk,rst,matrix_A[3345],matrix_B[145],mul_res1[3345]);
multi_7x28 multi_7x28_mod_3346(clk,rst,matrix_A[3346],matrix_B[146],mul_res1[3346]);
multi_7x28 multi_7x28_mod_3347(clk,rst,matrix_A[3347],matrix_B[147],mul_res1[3347]);
multi_7x28 multi_7x28_mod_3348(clk,rst,matrix_A[3348],matrix_B[148],mul_res1[3348]);
multi_7x28 multi_7x28_mod_3349(clk,rst,matrix_A[3349],matrix_B[149],mul_res1[3349]);
multi_7x28 multi_7x28_mod_3350(clk,rst,matrix_A[3350],matrix_B[150],mul_res1[3350]);
multi_7x28 multi_7x28_mod_3351(clk,rst,matrix_A[3351],matrix_B[151],mul_res1[3351]);
multi_7x28 multi_7x28_mod_3352(clk,rst,matrix_A[3352],matrix_B[152],mul_res1[3352]);
multi_7x28 multi_7x28_mod_3353(clk,rst,matrix_A[3353],matrix_B[153],mul_res1[3353]);
multi_7x28 multi_7x28_mod_3354(clk,rst,matrix_A[3354],matrix_B[154],mul_res1[3354]);
multi_7x28 multi_7x28_mod_3355(clk,rst,matrix_A[3355],matrix_B[155],mul_res1[3355]);
multi_7x28 multi_7x28_mod_3356(clk,rst,matrix_A[3356],matrix_B[156],mul_res1[3356]);
multi_7x28 multi_7x28_mod_3357(clk,rst,matrix_A[3357],matrix_B[157],mul_res1[3357]);
multi_7x28 multi_7x28_mod_3358(clk,rst,matrix_A[3358],matrix_B[158],mul_res1[3358]);
multi_7x28 multi_7x28_mod_3359(clk,rst,matrix_A[3359],matrix_B[159],mul_res1[3359]);
multi_7x28 multi_7x28_mod_3360(clk,rst,matrix_A[3360],matrix_B[160],mul_res1[3360]);
multi_7x28 multi_7x28_mod_3361(clk,rst,matrix_A[3361],matrix_B[161],mul_res1[3361]);
multi_7x28 multi_7x28_mod_3362(clk,rst,matrix_A[3362],matrix_B[162],mul_res1[3362]);
multi_7x28 multi_7x28_mod_3363(clk,rst,matrix_A[3363],matrix_B[163],mul_res1[3363]);
multi_7x28 multi_7x28_mod_3364(clk,rst,matrix_A[3364],matrix_B[164],mul_res1[3364]);
multi_7x28 multi_7x28_mod_3365(clk,rst,matrix_A[3365],matrix_B[165],mul_res1[3365]);
multi_7x28 multi_7x28_mod_3366(clk,rst,matrix_A[3366],matrix_B[166],mul_res1[3366]);
multi_7x28 multi_7x28_mod_3367(clk,rst,matrix_A[3367],matrix_B[167],mul_res1[3367]);
multi_7x28 multi_7x28_mod_3368(clk,rst,matrix_A[3368],matrix_B[168],mul_res1[3368]);
multi_7x28 multi_7x28_mod_3369(clk,rst,matrix_A[3369],matrix_B[169],mul_res1[3369]);
multi_7x28 multi_7x28_mod_3370(clk,rst,matrix_A[3370],matrix_B[170],mul_res1[3370]);
multi_7x28 multi_7x28_mod_3371(clk,rst,matrix_A[3371],matrix_B[171],mul_res1[3371]);
multi_7x28 multi_7x28_mod_3372(clk,rst,matrix_A[3372],matrix_B[172],mul_res1[3372]);
multi_7x28 multi_7x28_mod_3373(clk,rst,matrix_A[3373],matrix_B[173],mul_res1[3373]);
multi_7x28 multi_7x28_mod_3374(clk,rst,matrix_A[3374],matrix_B[174],mul_res1[3374]);
multi_7x28 multi_7x28_mod_3375(clk,rst,matrix_A[3375],matrix_B[175],mul_res1[3375]);
multi_7x28 multi_7x28_mod_3376(clk,rst,matrix_A[3376],matrix_B[176],mul_res1[3376]);
multi_7x28 multi_7x28_mod_3377(clk,rst,matrix_A[3377],matrix_B[177],mul_res1[3377]);
multi_7x28 multi_7x28_mod_3378(clk,rst,matrix_A[3378],matrix_B[178],mul_res1[3378]);
multi_7x28 multi_7x28_mod_3379(clk,rst,matrix_A[3379],matrix_B[179],mul_res1[3379]);
multi_7x28 multi_7x28_mod_3380(clk,rst,matrix_A[3380],matrix_B[180],mul_res1[3380]);
multi_7x28 multi_7x28_mod_3381(clk,rst,matrix_A[3381],matrix_B[181],mul_res1[3381]);
multi_7x28 multi_7x28_mod_3382(clk,rst,matrix_A[3382],matrix_B[182],mul_res1[3382]);
multi_7x28 multi_7x28_mod_3383(clk,rst,matrix_A[3383],matrix_B[183],mul_res1[3383]);
multi_7x28 multi_7x28_mod_3384(clk,rst,matrix_A[3384],matrix_B[184],mul_res1[3384]);
multi_7x28 multi_7x28_mod_3385(clk,rst,matrix_A[3385],matrix_B[185],mul_res1[3385]);
multi_7x28 multi_7x28_mod_3386(clk,rst,matrix_A[3386],matrix_B[186],mul_res1[3386]);
multi_7x28 multi_7x28_mod_3387(clk,rst,matrix_A[3387],matrix_B[187],mul_res1[3387]);
multi_7x28 multi_7x28_mod_3388(clk,rst,matrix_A[3388],matrix_B[188],mul_res1[3388]);
multi_7x28 multi_7x28_mod_3389(clk,rst,matrix_A[3389],matrix_B[189],mul_res1[3389]);
multi_7x28 multi_7x28_mod_3390(clk,rst,matrix_A[3390],matrix_B[190],mul_res1[3390]);
multi_7x28 multi_7x28_mod_3391(clk,rst,matrix_A[3391],matrix_B[191],mul_res1[3391]);
multi_7x28 multi_7x28_mod_3392(clk,rst,matrix_A[3392],matrix_B[192],mul_res1[3392]);
multi_7x28 multi_7x28_mod_3393(clk,rst,matrix_A[3393],matrix_B[193],mul_res1[3393]);
multi_7x28 multi_7x28_mod_3394(clk,rst,matrix_A[3394],matrix_B[194],mul_res1[3394]);
multi_7x28 multi_7x28_mod_3395(clk,rst,matrix_A[3395],matrix_B[195],mul_res1[3395]);
multi_7x28 multi_7x28_mod_3396(clk,rst,matrix_A[3396],matrix_B[196],mul_res1[3396]);
multi_7x28 multi_7x28_mod_3397(clk,rst,matrix_A[3397],matrix_B[197],mul_res1[3397]);
multi_7x28 multi_7x28_mod_3398(clk,rst,matrix_A[3398],matrix_B[198],mul_res1[3398]);
multi_7x28 multi_7x28_mod_3399(clk,rst,matrix_A[3399],matrix_B[199],mul_res1[3399]);
multi_7x28 multi_7x28_mod_3400(clk,rst,matrix_A[3400],matrix_B[0],mul_res1[3400]);
multi_7x28 multi_7x28_mod_3401(clk,rst,matrix_A[3401],matrix_B[1],mul_res1[3401]);
multi_7x28 multi_7x28_mod_3402(clk,rst,matrix_A[3402],matrix_B[2],mul_res1[3402]);
multi_7x28 multi_7x28_mod_3403(clk,rst,matrix_A[3403],matrix_B[3],mul_res1[3403]);
multi_7x28 multi_7x28_mod_3404(clk,rst,matrix_A[3404],matrix_B[4],mul_res1[3404]);
multi_7x28 multi_7x28_mod_3405(clk,rst,matrix_A[3405],matrix_B[5],mul_res1[3405]);
multi_7x28 multi_7x28_mod_3406(clk,rst,matrix_A[3406],matrix_B[6],mul_res1[3406]);
multi_7x28 multi_7x28_mod_3407(clk,rst,matrix_A[3407],matrix_B[7],mul_res1[3407]);
multi_7x28 multi_7x28_mod_3408(clk,rst,matrix_A[3408],matrix_B[8],mul_res1[3408]);
multi_7x28 multi_7x28_mod_3409(clk,rst,matrix_A[3409],matrix_B[9],mul_res1[3409]);
multi_7x28 multi_7x28_mod_3410(clk,rst,matrix_A[3410],matrix_B[10],mul_res1[3410]);
multi_7x28 multi_7x28_mod_3411(clk,rst,matrix_A[3411],matrix_B[11],mul_res1[3411]);
multi_7x28 multi_7x28_mod_3412(clk,rst,matrix_A[3412],matrix_B[12],mul_res1[3412]);
multi_7x28 multi_7x28_mod_3413(clk,rst,matrix_A[3413],matrix_B[13],mul_res1[3413]);
multi_7x28 multi_7x28_mod_3414(clk,rst,matrix_A[3414],matrix_B[14],mul_res1[3414]);
multi_7x28 multi_7x28_mod_3415(clk,rst,matrix_A[3415],matrix_B[15],mul_res1[3415]);
multi_7x28 multi_7x28_mod_3416(clk,rst,matrix_A[3416],matrix_B[16],mul_res1[3416]);
multi_7x28 multi_7x28_mod_3417(clk,rst,matrix_A[3417],matrix_B[17],mul_res1[3417]);
multi_7x28 multi_7x28_mod_3418(clk,rst,matrix_A[3418],matrix_B[18],mul_res1[3418]);
multi_7x28 multi_7x28_mod_3419(clk,rst,matrix_A[3419],matrix_B[19],mul_res1[3419]);
multi_7x28 multi_7x28_mod_3420(clk,rst,matrix_A[3420],matrix_B[20],mul_res1[3420]);
multi_7x28 multi_7x28_mod_3421(clk,rst,matrix_A[3421],matrix_B[21],mul_res1[3421]);
multi_7x28 multi_7x28_mod_3422(clk,rst,matrix_A[3422],matrix_B[22],mul_res1[3422]);
multi_7x28 multi_7x28_mod_3423(clk,rst,matrix_A[3423],matrix_B[23],mul_res1[3423]);
multi_7x28 multi_7x28_mod_3424(clk,rst,matrix_A[3424],matrix_B[24],mul_res1[3424]);
multi_7x28 multi_7x28_mod_3425(clk,rst,matrix_A[3425],matrix_B[25],mul_res1[3425]);
multi_7x28 multi_7x28_mod_3426(clk,rst,matrix_A[3426],matrix_B[26],mul_res1[3426]);
multi_7x28 multi_7x28_mod_3427(clk,rst,matrix_A[3427],matrix_B[27],mul_res1[3427]);
multi_7x28 multi_7x28_mod_3428(clk,rst,matrix_A[3428],matrix_B[28],mul_res1[3428]);
multi_7x28 multi_7x28_mod_3429(clk,rst,matrix_A[3429],matrix_B[29],mul_res1[3429]);
multi_7x28 multi_7x28_mod_3430(clk,rst,matrix_A[3430],matrix_B[30],mul_res1[3430]);
multi_7x28 multi_7x28_mod_3431(clk,rst,matrix_A[3431],matrix_B[31],mul_res1[3431]);
multi_7x28 multi_7x28_mod_3432(clk,rst,matrix_A[3432],matrix_B[32],mul_res1[3432]);
multi_7x28 multi_7x28_mod_3433(clk,rst,matrix_A[3433],matrix_B[33],mul_res1[3433]);
multi_7x28 multi_7x28_mod_3434(clk,rst,matrix_A[3434],matrix_B[34],mul_res1[3434]);
multi_7x28 multi_7x28_mod_3435(clk,rst,matrix_A[3435],matrix_B[35],mul_res1[3435]);
multi_7x28 multi_7x28_mod_3436(clk,rst,matrix_A[3436],matrix_B[36],mul_res1[3436]);
multi_7x28 multi_7x28_mod_3437(clk,rst,matrix_A[3437],matrix_B[37],mul_res1[3437]);
multi_7x28 multi_7x28_mod_3438(clk,rst,matrix_A[3438],matrix_B[38],mul_res1[3438]);
multi_7x28 multi_7x28_mod_3439(clk,rst,matrix_A[3439],matrix_B[39],mul_res1[3439]);
multi_7x28 multi_7x28_mod_3440(clk,rst,matrix_A[3440],matrix_B[40],mul_res1[3440]);
multi_7x28 multi_7x28_mod_3441(clk,rst,matrix_A[3441],matrix_B[41],mul_res1[3441]);
multi_7x28 multi_7x28_mod_3442(clk,rst,matrix_A[3442],matrix_B[42],mul_res1[3442]);
multi_7x28 multi_7x28_mod_3443(clk,rst,matrix_A[3443],matrix_B[43],mul_res1[3443]);
multi_7x28 multi_7x28_mod_3444(clk,rst,matrix_A[3444],matrix_B[44],mul_res1[3444]);
multi_7x28 multi_7x28_mod_3445(clk,rst,matrix_A[3445],matrix_B[45],mul_res1[3445]);
multi_7x28 multi_7x28_mod_3446(clk,rst,matrix_A[3446],matrix_B[46],mul_res1[3446]);
multi_7x28 multi_7x28_mod_3447(clk,rst,matrix_A[3447],matrix_B[47],mul_res1[3447]);
multi_7x28 multi_7x28_mod_3448(clk,rst,matrix_A[3448],matrix_B[48],mul_res1[3448]);
multi_7x28 multi_7x28_mod_3449(clk,rst,matrix_A[3449],matrix_B[49],mul_res1[3449]);
multi_7x28 multi_7x28_mod_3450(clk,rst,matrix_A[3450],matrix_B[50],mul_res1[3450]);
multi_7x28 multi_7x28_mod_3451(clk,rst,matrix_A[3451],matrix_B[51],mul_res1[3451]);
multi_7x28 multi_7x28_mod_3452(clk,rst,matrix_A[3452],matrix_B[52],mul_res1[3452]);
multi_7x28 multi_7x28_mod_3453(clk,rst,matrix_A[3453],matrix_B[53],mul_res1[3453]);
multi_7x28 multi_7x28_mod_3454(clk,rst,matrix_A[3454],matrix_B[54],mul_res1[3454]);
multi_7x28 multi_7x28_mod_3455(clk,rst,matrix_A[3455],matrix_B[55],mul_res1[3455]);
multi_7x28 multi_7x28_mod_3456(clk,rst,matrix_A[3456],matrix_B[56],mul_res1[3456]);
multi_7x28 multi_7x28_mod_3457(clk,rst,matrix_A[3457],matrix_B[57],mul_res1[3457]);
multi_7x28 multi_7x28_mod_3458(clk,rst,matrix_A[3458],matrix_B[58],mul_res1[3458]);
multi_7x28 multi_7x28_mod_3459(clk,rst,matrix_A[3459],matrix_B[59],mul_res1[3459]);
multi_7x28 multi_7x28_mod_3460(clk,rst,matrix_A[3460],matrix_B[60],mul_res1[3460]);
multi_7x28 multi_7x28_mod_3461(clk,rst,matrix_A[3461],matrix_B[61],mul_res1[3461]);
multi_7x28 multi_7x28_mod_3462(clk,rst,matrix_A[3462],matrix_B[62],mul_res1[3462]);
multi_7x28 multi_7x28_mod_3463(clk,rst,matrix_A[3463],matrix_B[63],mul_res1[3463]);
multi_7x28 multi_7x28_mod_3464(clk,rst,matrix_A[3464],matrix_B[64],mul_res1[3464]);
multi_7x28 multi_7x28_mod_3465(clk,rst,matrix_A[3465],matrix_B[65],mul_res1[3465]);
multi_7x28 multi_7x28_mod_3466(clk,rst,matrix_A[3466],matrix_B[66],mul_res1[3466]);
multi_7x28 multi_7x28_mod_3467(clk,rst,matrix_A[3467],matrix_B[67],mul_res1[3467]);
multi_7x28 multi_7x28_mod_3468(clk,rst,matrix_A[3468],matrix_B[68],mul_res1[3468]);
multi_7x28 multi_7x28_mod_3469(clk,rst,matrix_A[3469],matrix_B[69],mul_res1[3469]);
multi_7x28 multi_7x28_mod_3470(clk,rst,matrix_A[3470],matrix_B[70],mul_res1[3470]);
multi_7x28 multi_7x28_mod_3471(clk,rst,matrix_A[3471],matrix_B[71],mul_res1[3471]);
multi_7x28 multi_7x28_mod_3472(clk,rst,matrix_A[3472],matrix_B[72],mul_res1[3472]);
multi_7x28 multi_7x28_mod_3473(clk,rst,matrix_A[3473],matrix_B[73],mul_res1[3473]);
multi_7x28 multi_7x28_mod_3474(clk,rst,matrix_A[3474],matrix_B[74],mul_res1[3474]);
multi_7x28 multi_7x28_mod_3475(clk,rst,matrix_A[3475],matrix_B[75],mul_res1[3475]);
multi_7x28 multi_7x28_mod_3476(clk,rst,matrix_A[3476],matrix_B[76],mul_res1[3476]);
multi_7x28 multi_7x28_mod_3477(clk,rst,matrix_A[3477],matrix_B[77],mul_res1[3477]);
multi_7x28 multi_7x28_mod_3478(clk,rst,matrix_A[3478],matrix_B[78],mul_res1[3478]);
multi_7x28 multi_7x28_mod_3479(clk,rst,matrix_A[3479],matrix_B[79],mul_res1[3479]);
multi_7x28 multi_7x28_mod_3480(clk,rst,matrix_A[3480],matrix_B[80],mul_res1[3480]);
multi_7x28 multi_7x28_mod_3481(clk,rst,matrix_A[3481],matrix_B[81],mul_res1[3481]);
multi_7x28 multi_7x28_mod_3482(clk,rst,matrix_A[3482],matrix_B[82],mul_res1[3482]);
multi_7x28 multi_7x28_mod_3483(clk,rst,matrix_A[3483],matrix_B[83],mul_res1[3483]);
multi_7x28 multi_7x28_mod_3484(clk,rst,matrix_A[3484],matrix_B[84],mul_res1[3484]);
multi_7x28 multi_7x28_mod_3485(clk,rst,matrix_A[3485],matrix_B[85],mul_res1[3485]);
multi_7x28 multi_7x28_mod_3486(clk,rst,matrix_A[3486],matrix_B[86],mul_res1[3486]);
multi_7x28 multi_7x28_mod_3487(clk,rst,matrix_A[3487],matrix_B[87],mul_res1[3487]);
multi_7x28 multi_7x28_mod_3488(clk,rst,matrix_A[3488],matrix_B[88],mul_res1[3488]);
multi_7x28 multi_7x28_mod_3489(clk,rst,matrix_A[3489],matrix_B[89],mul_res1[3489]);
multi_7x28 multi_7x28_mod_3490(clk,rst,matrix_A[3490],matrix_B[90],mul_res1[3490]);
multi_7x28 multi_7x28_mod_3491(clk,rst,matrix_A[3491],matrix_B[91],mul_res1[3491]);
multi_7x28 multi_7x28_mod_3492(clk,rst,matrix_A[3492],matrix_B[92],mul_res1[3492]);
multi_7x28 multi_7x28_mod_3493(clk,rst,matrix_A[3493],matrix_B[93],mul_res1[3493]);
multi_7x28 multi_7x28_mod_3494(clk,rst,matrix_A[3494],matrix_B[94],mul_res1[3494]);
multi_7x28 multi_7x28_mod_3495(clk,rst,matrix_A[3495],matrix_B[95],mul_res1[3495]);
multi_7x28 multi_7x28_mod_3496(clk,rst,matrix_A[3496],matrix_B[96],mul_res1[3496]);
multi_7x28 multi_7x28_mod_3497(clk,rst,matrix_A[3497],matrix_B[97],mul_res1[3497]);
multi_7x28 multi_7x28_mod_3498(clk,rst,matrix_A[3498],matrix_B[98],mul_res1[3498]);
multi_7x28 multi_7x28_mod_3499(clk,rst,matrix_A[3499],matrix_B[99],mul_res1[3499]);
multi_7x28 multi_7x28_mod_3500(clk,rst,matrix_A[3500],matrix_B[100],mul_res1[3500]);
multi_7x28 multi_7x28_mod_3501(clk,rst,matrix_A[3501],matrix_B[101],mul_res1[3501]);
multi_7x28 multi_7x28_mod_3502(clk,rst,matrix_A[3502],matrix_B[102],mul_res1[3502]);
multi_7x28 multi_7x28_mod_3503(clk,rst,matrix_A[3503],matrix_B[103],mul_res1[3503]);
multi_7x28 multi_7x28_mod_3504(clk,rst,matrix_A[3504],matrix_B[104],mul_res1[3504]);
multi_7x28 multi_7x28_mod_3505(clk,rst,matrix_A[3505],matrix_B[105],mul_res1[3505]);
multi_7x28 multi_7x28_mod_3506(clk,rst,matrix_A[3506],matrix_B[106],mul_res1[3506]);
multi_7x28 multi_7x28_mod_3507(clk,rst,matrix_A[3507],matrix_B[107],mul_res1[3507]);
multi_7x28 multi_7x28_mod_3508(clk,rst,matrix_A[3508],matrix_B[108],mul_res1[3508]);
multi_7x28 multi_7x28_mod_3509(clk,rst,matrix_A[3509],matrix_B[109],mul_res1[3509]);
multi_7x28 multi_7x28_mod_3510(clk,rst,matrix_A[3510],matrix_B[110],mul_res1[3510]);
multi_7x28 multi_7x28_mod_3511(clk,rst,matrix_A[3511],matrix_B[111],mul_res1[3511]);
multi_7x28 multi_7x28_mod_3512(clk,rst,matrix_A[3512],matrix_B[112],mul_res1[3512]);
multi_7x28 multi_7x28_mod_3513(clk,rst,matrix_A[3513],matrix_B[113],mul_res1[3513]);
multi_7x28 multi_7x28_mod_3514(clk,rst,matrix_A[3514],matrix_B[114],mul_res1[3514]);
multi_7x28 multi_7x28_mod_3515(clk,rst,matrix_A[3515],matrix_B[115],mul_res1[3515]);
multi_7x28 multi_7x28_mod_3516(clk,rst,matrix_A[3516],matrix_B[116],mul_res1[3516]);
multi_7x28 multi_7x28_mod_3517(clk,rst,matrix_A[3517],matrix_B[117],mul_res1[3517]);
multi_7x28 multi_7x28_mod_3518(clk,rst,matrix_A[3518],matrix_B[118],mul_res1[3518]);
multi_7x28 multi_7x28_mod_3519(clk,rst,matrix_A[3519],matrix_B[119],mul_res1[3519]);
multi_7x28 multi_7x28_mod_3520(clk,rst,matrix_A[3520],matrix_B[120],mul_res1[3520]);
multi_7x28 multi_7x28_mod_3521(clk,rst,matrix_A[3521],matrix_B[121],mul_res1[3521]);
multi_7x28 multi_7x28_mod_3522(clk,rst,matrix_A[3522],matrix_B[122],mul_res1[3522]);
multi_7x28 multi_7x28_mod_3523(clk,rst,matrix_A[3523],matrix_B[123],mul_res1[3523]);
multi_7x28 multi_7x28_mod_3524(clk,rst,matrix_A[3524],matrix_B[124],mul_res1[3524]);
multi_7x28 multi_7x28_mod_3525(clk,rst,matrix_A[3525],matrix_B[125],mul_res1[3525]);
multi_7x28 multi_7x28_mod_3526(clk,rst,matrix_A[3526],matrix_B[126],mul_res1[3526]);
multi_7x28 multi_7x28_mod_3527(clk,rst,matrix_A[3527],matrix_B[127],mul_res1[3527]);
multi_7x28 multi_7x28_mod_3528(clk,rst,matrix_A[3528],matrix_B[128],mul_res1[3528]);
multi_7x28 multi_7x28_mod_3529(clk,rst,matrix_A[3529],matrix_B[129],mul_res1[3529]);
multi_7x28 multi_7x28_mod_3530(clk,rst,matrix_A[3530],matrix_B[130],mul_res1[3530]);
multi_7x28 multi_7x28_mod_3531(clk,rst,matrix_A[3531],matrix_B[131],mul_res1[3531]);
multi_7x28 multi_7x28_mod_3532(clk,rst,matrix_A[3532],matrix_B[132],mul_res1[3532]);
multi_7x28 multi_7x28_mod_3533(clk,rst,matrix_A[3533],matrix_B[133],mul_res1[3533]);
multi_7x28 multi_7x28_mod_3534(clk,rst,matrix_A[3534],matrix_B[134],mul_res1[3534]);
multi_7x28 multi_7x28_mod_3535(clk,rst,matrix_A[3535],matrix_B[135],mul_res1[3535]);
multi_7x28 multi_7x28_mod_3536(clk,rst,matrix_A[3536],matrix_B[136],mul_res1[3536]);
multi_7x28 multi_7x28_mod_3537(clk,rst,matrix_A[3537],matrix_B[137],mul_res1[3537]);
multi_7x28 multi_7x28_mod_3538(clk,rst,matrix_A[3538],matrix_B[138],mul_res1[3538]);
multi_7x28 multi_7x28_mod_3539(clk,rst,matrix_A[3539],matrix_B[139],mul_res1[3539]);
multi_7x28 multi_7x28_mod_3540(clk,rst,matrix_A[3540],matrix_B[140],mul_res1[3540]);
multi_7x28 multi_7x28_mod_3541(clk,rst,matrix_A[3541],matrix_B[141],mul_res1[3541]);
multi_7x28 multi_7x28_mod_3542(clk,rst,matrix_A[3542],matrix_B[142],mul_res1[3542]);
multi_7x28 multi_7x28_mod_3543(clk,rst,matrix_A[3543],matrix_B[143],mul_res1[3543]);
multi_7x28 multi_7x28_mod_3544(clk,rst,matrix_A[3544],matrix_B[144],mul_res1[3544]);
multi_7x28 multi_7x28_mod_3545(clk,rst,matrix_A[3545],matrix_B[145],mul_res1[3545]);
multi_7x28 multi_7x28_mod_3546(clk,rst,matrix_A[3546],matrix_B[146],mul_res1[3546]);
multi_7x28 multi_7x28_mod_3547(clk,rst,matrix_A[3547],matrix_B[147],mul_res1[3547]);
multi_7x28 multi_7x28_mod_3548(clk,rst,matrix_A[3548],matrix_B[148],mul_res1[3548]);
multi_7x28 multi_7x28_mod_3549(clk,rst,matrix_A[3549],matrix_B[149],mul_res1[3549]);
multi_7x28 multi_7x28_mod_3550(clk,rst,matrix_A[3550],matrix_B[150],mul_res1[3550]);
multi_7x28 multi_7x28_mod_3551(clk,rst,matrix_A[3551],matrix_B[151],mul_res1[3551]);
multi_7x28 multi_7x28_mod_3552(clk,rst,matrix_A[3552],matrix_B[152],mul_res1[3552]);
multi_7x28 multi_7x28_mod_3553(clk,rst,matrix_A[3553],matrix_B[153],mul_res1[3553]);
multi_7x28 multi_7x28_mod_3554(clk,rst,matrix_A[3554],matrix_B[154],mul_res1[3554]);
multi_7x28 multi_7x28_mod_3555(clk,rst,matrix_A[3555],matrix_B[155],mul_res1[3555]);
multi_7x28 multi_7x28_mod_3556(clk,rst,matrix_A[3556],matrix_B[156],mul_res1[3556]);
multi_7x28 multi_7x28_mod_3557(clk,rst,matrix_A[3557],matrix_B[157],mul_res1[3557]);
multi_7x28 multi_7x28_mod_3558(clk,rst,matrix_A[3558],matrix_B[158],mul_res1[3558]);
multi_7x28 multi_7x28_mod_3559(clk,rst,matrix_A[3559],matrix_B[159],mul_res1[3559]);
multi_7x28 multi_7x28_mod_3560(clk,rst,matrix_A[3560],matrix_B[160],mul_res1[3560]);
multi_7x28 multi_7x28_mod_3561(clk,rst,matrix_A[3561],matrix_B[161],mul_res1[3561]);
multi_7x28 multi_7x28_mod_3562(clk,rst,matrix_A[3562],matrix_B[162],mul_res1[3562]);
multi_7x28 multi_7x28_mod_3563(clk,rst,matrix_A[3563],matrix_B[163],mul_res1[3563]);
multi_7x28 multi_7x28_mod_3564(clk,rst,matrix_A[3564],matrix_B[164],mul_res1[3564]);
multi_7x28 multi_7x28_mod_3565(clk,rst,matrix_A[3565],matrix_B[165],mul_res1[3565]);
multi_7x28 multi_7x28_mod_3566(clk,rst,matrix_A[3566],matrix_B[166],mul_res1[3566]);
multi_7x28 multi_7x28_mod_3567(clk,rst,matrix_A[3567],matrix_B[167],mul_res1[3567]);
multi_7x28 multi_7x28_mod_3568(clk,rst,matrix_A[3568],matrix_B[168],mul_res1[3568]);
multi_7x28 multi_7x28_mod_3569(clk,rst,matrix_A[3569],matrix_B[169],mul_res1[3569]);
multi_7x28 multi_7x28_mod_3570(clk,rst,matrix_A[3570],matrix_B[170],mul_res1[3570]);
multi_7x28 multi_7x28_mod_3571(clk,rst,matrix_A[3571],matrix_B[171],mul_res1[3571]);
multi_7x28 multi_7x28_mod_3572(clk,rst,matrix_A[3572],matrix_B[172],mul_res1[3572]);
multi_7x28 multi_7x28_mod_3573(clk,rst,matrix_A[3573],matrix_B[173],mul_res1[3573]);
multi_7x28 multi_7x28_mod_3574(clk,rst,matrix_A[3574],matrix_B[174],mul_res1[3574]);
multi_7x28 multi_7x28_mod_3575(clk,rst,matrix_A[3575],matrix_B[175],mul_res1[3575]);
multi_7x28 multi_7x28_mod_3576(clk,rst,matrix_A[3576],matrix_B[176],mul_res1[3576]);
multi_7x28 multi_7x28_mod_3577(clk,rst,matrix_A[3577],matrix_B[177],mul_res1[3577]);
multi_7x28 multi_7x28_mod_3578(clk,rst,matrix_A[3578],matrix_B[178],mul_res1[3578]);
multi_7x28 multi_7x28_mod_3579(clk,rst,matrix_A[3579],matrix_B[179],mul_res1[3579]);
multi_7x28 multi_7x28_mod_3580(clk,rst,matrix_A[3580],matrix_B[180],mul_res1[3580]);
multi_7x28 multi_7x28_mod_3581(clk,rst,matrix_A[3581],matrix_B[181],mul_res1[3581]);
multi_7x28 multi_7x28_mod_3582(clk,rst,matrix_A[3582],matrix_B[182],mul_res1[3582]);
multi_7x28 multi_7x28_mod_3583(clk,rst,matrix_A[3583],matrix_B[183],mul_res1[3583]);
multi_7x28 multi_7x28_mod_3584(clk,rst,matrix_A[3584],matrix_B[184],mul_res1[3584]);
multi_7x28 multi_7x28_mod_3585(clk,rst,matrix_A[3585],matrix_B[185],mul_res1[3585]);
multi_7x28 multi_7x28_mod_3586(clk,rst,matrix_A[3586],matrix_B[186],mul_res1[3586]);
multi_7x28 multi_7x28_mod_3587(clk,rst,matrix_A[3587],matrix_B[187],mul_res1[3587]);
multi_7x28 multi_7x28_mod_3588(clk,rst,matrix_A[3588],matrix_B[188],mul_res1[3588]);
multi_7x28 multi_7x28_mod_3589(clk,rst,matrix_A[3589],matrix_B[189],mul_res1[3589]);
multi_7x28 multi_7x28_mod_3590(clk,rst,matrix_A[3590],matrix_B[190],mul_res1[3590]);
multi_7x28 multi_7x28_mod_3591(clk,rst,matrix_A[3591],matrix_B[191],mul_res1[3591]);
multi_7x28 multi_7x28_mod_3592(clk,rst,matrix_A[3592],matrix_B[192],mul_res1[3592]);
multi_7x28 multi_7x28_mod_3593(clk,rst,matrix_A[3593],matrix_B[193],mul_res1[3593]);
multi_7x28 multi_7x28_mod_3594(clk,rst,matrix_A[3594],matrix_B[194],mul_res1[3594]);
multi_7x28 multi_7x28_mod_3595(clk,rst,matrix_A[3595],matrix_B[195],mul_res1[3595]);
multi_7x28 multi_7x28_mod_3596(clk,rst,matrix_A[3596],matrix_B[196],mul_res1[3596]);
multi_7x28 multi_7x28_mod_3597(clk,rst,matrix_A[3597],matrix_B[197],mul_res1[3597]);
multi_7x28 multi_7x28_mod_3598(clk,rst,matrix_A[3598],matrix_B[198],mul_res1[3598]);
multi_7x28 multi_7x28_mod_3599(clk,rst,matrix_A[3599],matrix_B[199],mul_res1[3599]);
multi_7x28 multi_7x28_mod_3600(clk,rst,matrix_A[3600],matrix_B[0],mul_res1[3600]);
multi_7x28 multi_7x28_mod_3601(clk,rst,matrix_A[3601],matrix_B[1],mul_res1[3601]);
multi_7x28 multi_7x28_mod_3602(clk,rst,matrix_A[3602],matrix_B[2],mul_res1[3602]);
multi_7x28 multi_7x28_mod_3603(clk,rst,matrix_A[3603],matrix_B[3],mul_res1[3603]);
multi_7x28 multi_7x28_mod_3604(clk,rst,matrix_A[3604],matrix_B[4],mul_res1[3604]);
multi_7x28 multi_7x28_mod_3605(clk,rst,matrix_A[3605],matrix_B[5],mul_res1[3605]);
multi_7x28 multi_7x28_mod_3606(clk,rst,matrix_A[3606],matrix_B[6],mul_res1[3606]);
multi_7x28 multi_7x28_mod_3607(clk,rst,matrix_A[3607],matrix_B[7],mul_res1[3607]);
multi_7x28 multi_7x28_mod_3608(clk,rst,matrix_A[3608],matrix_B[8],mul_res1[3608]);
multi_7x28 multi_7x28_mod_3609(clk,rst,matrix_A[3609],matrix_B[9],mul_res1[3609]);
multi_7x28 multi_7x28_mod_3610(clk,rst,matrix_A[3610],matrix_B[10],mul_res1[3610]);
multi_7x28 multi_7x28_mod_3611(clk,rst,matrix_A[3611],matrix_B[11],mul_res1[3611]);
multi_7x28 multi_7x28_mod_3612(clk,rst,matrix_A[3612],matrix_B[12],mul_res1[3612]);
multi_7x28 multi_7x28_mod_3613(clk,rst,matrix_A[3613],matrix_B[13],mul_res1[3613]);
multi_7x28 multi_7x28_mod_3614(clk,rst,matrix_A[3614],matrix_B[14],mul_res1[3614]);
multi_7x28 multi_7x28_mod_3615(clk,rst,matrix_A[3615],matrix_B[15],mul_res1[3615]);
multi_7x28 multi_7x28_mod_3616(clk,rst,matrix_A[3616],matrix_B[16],mul_res1[3616]);
multi_7x28 multi_7x28_mod_3617(clk,rst,matrix_A[3617],matrix_B[17],mul_res1[3617]);
multi_7x28 multi_7x28_mod_3618(clk,rst,matrix_A[3618],matrix_B[18],mul_res1[3618]);
multi_7x28 multi_7x28_mod_3619(clk,rst,matrix_A[3619],matrix_B[19],mul_res1[3619]);
multi_7x28 multi_7x28_mod_3620(clk,rst,matrix_A[3620],matrix_B[20],mul_res1[3620]);
multi_7x28 multi_7x28_mod_3621(clk,rst,matrix_A[3621],matrix_B[21],mul_res1[3621]);
multi_7x28 multi_7x28_mod_3622(clk,rst,matrix_A[3622],matrix_B[22],mul_res1[3622]);
multi_7x28 multi_7x28_mod_3623(clk,rst,matrix_A[3623],matrix_B[23],mul_res1[3623]);
multi_7x28 multi_7x28_mod_3624(clk,rst,matrix_A[3624],matrix_B[24],mul_res1[3624]);
multi_7x28 multi_7x28_mod_3625(clk,rst,matrix_A[3625],matrix_B[25],mul_res1[3625]);
multi_7x28 multi_7x28_mod_3626(clk,rst,matrix_A[3626],matrix_B[26],mul_res1[3626]);
multi_7x28 multi_7x28_mod_3627(clk,rst,matrix_A[3627],matrix_B[27],mul_res1[3627]);
multi_7x28 multi_7x28_mod_3628(clk,rst,matrix_A[3628],matrix_B[28],mul_res1[3628]);
multi_7x28 multi_7x28_mod_3629(clk,rst,matrix_A[3629],matrix_B[29],mul_res1[3629]);
multi_7x28 multi_7x28_mod_3630(clk,rst,matrix_A[3630],matrix_B[30],mul_res1[3630]);
multi_7x28 multi_7x28_mod_3631(clk,rst,matrix_A[3631],matrix_B[31],mul_res1[3631]);
multi_7x28 multi_7x28_mod_3632(clk,rst,matrix_A[3632],matrix_B[32],mul_res1[3632]);
multi_7x28 multi_7x28_mod_3633(clk,rst,matrix_A[3633],matrix_B[33],mul_res1[3633]);
multi_7x28 multi_7x28_mod_3634(clk,rst,matrix_A[3634],matrix_B[34],mul_res1[3634]);
multi_7x28 multi_7x28_mod_3635(clk,rst,matrix_A[3635],matrix_B[35],mul_res1[3635]);
multi_7x28 multi_7x28_mod_3636(clk,rst,matrix_A[3636],matrix_B[36],mul_res1[3636]);
multi_7x28 multi_7x28_mod_3637(clk,rst,matrix_A[3637],matrix_B[37],mul_res1[3637]);
multi_7x28 multi_7x28_mod_3638(clk,rst,matrix_A[3638],matrix_B[38],mul_res1[3638]);
multi_7x28 multi_7x28_mod_3639(clk,rst,matrix_A[3639],matrix_B[39],mul_res1[3639]);
multi_7x28 multi_7x28_mod_3640(clk,rst,matrix_A[3640],matrix_B[40],mul_res1[3640]);
multi_7x28 multi_7x28_mod_3641(clk,rst,matrix_A[3641],matrix_B[41],mul_res1[3641]);
multi_7x28 multi_7x28_mod_3642(clk,rst,matrix_A[3642],matrix_B[42],mul_res1[3642]);
multi_7x28 multi_7x28_mod_3643(clk,rst,matrix_A[3643],matrix_B[43],mul_res1[3643]);
multi_7x28 multi_7x28_mod_3644(clk,rst,matrix_A[3644],matrix_B[44],mul_res1[3644]);
multi_7x28 multi_7x28_mod_3645(clk,rst,matrix_A[3645],matrix_B[45],mul_res1[3645]);
multi_7x28 multi_7x28_mod_3646(clk,rst,matrix_A[3646],matrix_B[46],mul_res1[3646]);
multi_7x28 multi_7x28_mod_3647(clk,rst,matrix_A[3647],matrix_B[47],mul_res1[3647]);
multi_7x28 multi_7x28_mod_3648(clk,rst,matrix_A[3648],matrix_B[48],mul_res1[3648]);
multi_7x28 multi_7x28_mod_3649(clk,rst,matrix_A[3649],matrix_B[49],mul_res1[3649]);
multi_7x28 multi_7x28_mod_3650(clk,rst,matrix_A[3650],matrix_B[50],mul_res1[3650]);
multi_7x28 multi_7x28_mod_3651(clk,rst,matrix_A[3651],matrix_B[51],mul_res1[3651]);
multi_7x28 multi_7x28_mod_3652(clk,rst,matrix_A[3652],matrix_B[52],mul_res1[3652]);
multi_7x28 multi_7x28_mod_3653(clk,rst,matrix_A[3653],matrix_B[53],mul_res1[3653]);
multi_7x28 multi_7x28_mod_3654(clk,rst,matrix_A[3654],matrix_B[54],mul_res1[3654]);
multi_7x28 multi_7x28_mod_3655(clk,rst,matrix_A[3655],matrix_B[55],mul_res1[3655]);
multi_7x28 multi_7x28_mod_3656(clk,rst,matrix_A[3656],matrix_B[56],mul_res1[3656]);
multi_7x28 multi_7x28_mod_3657(clk,rst,matrix_A[3657],matrix_B[57],mul_res1[3657]);
multi_7x28 multi_7x28_mod_3658(clk,rst,matrix_A[3658],matrix_B[58],mul_res1[3658]);
multi_7x28 multi_7x28_mod_3659(clk,rst,matrix_A[3659],matrix_B[59],mul_res1[3659]);
multi_7x28 multi_7x28_mod_3660(clk,rst,matrix_A[3660],matrix_B[60],mul_res1[3660]);
multi_7x28 multi_7x28_mod_3661(clk,rst,matrix_A[3661],matrix_B[61],mul_res1[3661]);
multi_7x28 multi_7x28_mod_3662(clk,rst,matrix_A[3662],matrix_B[62],mul_res1[3662]);
multi_7x28 multi_7x28_mod_3663(clk,rst,matrix_A[3663],matrix_B[63],mul_res1[3663]);
multi_7x28 multi_7x28_mod_3664(clk,rst,matrix_A[3664],matrix_B[64],mul_res1[3664]);
multi_7x28 multi_7x28_mod_3665(clk,rst,matrix_A[3665],matrix_B[65],mul_res1[3665]);
multi_7x28 multi_7x28_mod_3666(clk,rst,matrix_A[3666],matrix_B[66],mul_res1[3666]);
multi_7x28 multi_7x28_mod_3667(clk,rst,matrix_A[3667],matrix_B[67],mul_res1[3667]);
multi_7x28 multi_7x28_mod_3668(clk,rst,matrix_A[3668],matrix_B[68],mul_res1[3668]);
multi_7x28 multi_7x28_mod_3669(clk,rst,matrix_A[3669],matrix_B[69],mul_res1[3669]);
multi_7x28 multi_7x28_mod_3670(clk,rst,matrix_A[3670],matrix_B[70],mul_res1[3670]);
multi_7x28 multi_7x28_mod_3671(clk,rst,matrix_A[3671],matrix_B[71],mul_res1[3671]);
multi_7x28 multi_7x28_mod_3672(clk,rst,matrix_A[3672],matrix_B[72],mul_res1[3672]);
multi_7x28 multi_7x28_mod_3673(clk,rst,matrix_A[3673],matrix_B[73],mul_res1[3673]);
multi_7x28 multi_7x28_mod_3674(clk,rst,matrix_A[3674],matrix_B[74],mul_res1[3674]);
multi_7x28 multi_7x28_mod_3675(clk,rst,matrix_A[3675],matrix_B[75],mul_res1[3675]);
multi_7x28 multi_7x28_mod_3676(clk,rst,matrix_A[3676],matrix_B[76],mul_res1[3676]);
multi_7x28 multi_7x28_mod_3677(clk,rst,matrix_A[3677],matrix_B[77],mul_res1[3677]);
multi_7x28 multi_7x28_mod_3678(clk,rst,matrix_A[3678],matrix_B[78],mul_res1[3678]);
multi_7x28 multi_7x28_mod_3679(clk,rst,matrix_A[3679],matrix_B[79],mul_res1[3679]);
multi_7x28 multi_7x28_mod_3680(clk,rst,matrix_A[3680],matrix_B[80],mul_res1[3680]);
multi_7x28 multi_7x28_mod_3681(clk,rst,matrix_A[3681],matrix_B[81],mul_res1[3681]);
multi_7x28 multi_7x28_mod_3682(clk,rst,matrix_A[3682],matrix_B[82],mul_res1[3682]);
multi_7x28 multi_7x28_mod_3683(clk,rst,matrix_A[3683],matrix_B[83],mul_res1[3683]);
multi_7x28 multi_7x28_mod_3684(clk,rst,matrix_A[3684],matrix_B[84],mul_res1[3684]);
multi_7x28 multi_7x28_mod_3685(clk,rst,matrix_A[3685],matrix_B[85],mul_res1[3685]);
multi_7x28 multi_7x28_mod_3686(clk,rst,matrix_A[3686],matrix_B[86],mul_res1[3686]);
multi_7x28 multi_7x28_mod_3687(clk,rst,matrix_A[3687],matrix_B[87],mul_res1[3687]);
multi_7x28 multi_7x28_mod_3688(clk,rst,matrix_A[3688],matrix_B[88],mul_res1[3688]);
multi_7x28 multi_7x28_mod_3689(clk,rst,matrix_A[3689],matrix_B[89],mul_res1[3689]);
multi_7x28 multi_7x28_mod_3690(clk,rst,matrix_A[3690],matrix_B[90],mul_res1[3690]);
multi_7x28 multi_7x28_mod_3691(clk,rst,matrix_A[3691],matrix_B[91],mul_res1[3691]);
multi_7x28 multi_7x28_mod_3692(clk,rst,matrix_A[3692],matrix_B[92],mul_res1[3692]);
multi_7x28 multi_7x28_mod_3693(clk,rst,matrix_A[3693],matrix_B[93],mul_res1[3693]);
multi_7x28 multi_7x28_mod_3694(clk,rst,matrix_A[3694],matrix_B[94],mul_res1[3694]);
multi_7x28 multi_7x28_mod_3695(clk,rst,matrix_A[3695],matrix_B[95],mul_res1[3695]);
multi_7x28 multi_7x28_mod_3696(clk,rst,matrix_A[3696],matrix_B[96],mul_res1[3696]);
multi_7x28 multi_7x28_mod_3697(clk,rst,matrix_A[3697],matrix_B[97],mul_res1[3697]);
multi_7x28 multi_7x28_mod_3698(clk,rst,matrix_A[3698],matrix_B[98],mul_res1[3698]);
multi_7x28 multi_7x28_mod_3699(clk,rst,matrix_A[3699],matrix_B[99],mul_res1[3699]);
multi_7x28 multi_7x28_mod_3700(clk,rst,matrix_A[3700],matrix_B[100],mul_res1[3700]);
multi_7x28 multi_7x28_mod_3701(clk,rst,matrix_A[3701],matrix_B[101],mul_res1[3701]);
multi_7x28 multi_7x28_mod_3702(clk,rst,matrix_A[3702],matrix_B[102],mul_res1[3702]);
multi_7x28 multi_7x28_mod_3703(clk,rst,matrix_A[3703],matrix_B[103],mul_res1[3703]);
multi_7x28 multi_7x28_mod_3704(clk,rst,matrix_A[3704],matrix_B[104],mul_res1[3704]);
multi_7x28 multi_7x28_mod_3705(clk,rst,matrix_A[3705],matrix_B[105],mul_res1[3705]);
multi_7x28 multi_7x28_mod_3706(clk,rst,matrix_A[3706],matrix_B[106],mul_res1[3706]);
multi_7x28 multi_7x28_mod_3707(clk,rst,matrix_A[3707],matrix_B[107],mul_res1[3707]);
multi_7x28 multi_7x28_mod_3708(clk,rst,matrix_A[3708],matrix_B[108],mul_res1[3708]);
multi_7x28 multi_7x28_mod_3709(clk,rst,matrix_A[3709],matrix_B[109],mul_res1[3709]);
multi_7x28 multi_7x28_mod_3710(clk,rst,matrix_A[3710],matrix_B[110],mul_res1[3710]);
multi_7x28 multi_7x28_mod_3711(clk,rst,matrix_A[3711],matrix_B[111],mul_res1[3711]);
multi_7x28 multi_7x28_mod_3712(clk,rst,matrix_A[3712],matrix_B[112],mul_res1[3712]);
multi_7x28 multi_7x28_mod_3713(clk,rst,matrix_A[3713],matrix_B[113],mul_res1[3713]);
multi_7x28 multi_7x28_mod_3714(clk,rst,matrix_A[3714],matrix_B[114],mul_res1[3714]);
multi_7x28 multi_7x28_mod_3715(clk,rst,matrix_A[3715],matrix_B[115],mul_res1[3715]);
multi_7x28 multi_7x28_mod_3716(clk,rst,matrix_A[3716],matrix_B[116],mul_res1[3716]);
multi_7x28 multi_7x28_mod_3717(clk,rst,matrix_A[3717],matrix_B[117],mul_res1[3717]);
multi_7x28 multi_7x28_mod_3718(clk,rst,matrix_A[3718],matrix_B[118],mul_res1[3718]);
multi_7x28 multi_7x28_mod_3719(clk,rst,matrix_A[3719],matrix_B[119],mul_res1[3719]);
multi_7x28 multi_7x28_mod_3720(clk,rst,matrix_A[3720],matrix_B[120],mul_res1[3720]);
multi_7x28 multi_7x28_mod_3721(clk,rst,matrix_A[3721],matrix_B[121],mul_res1[3721]);
multi_7x28 multi_7x28_mod_3722(clk,rst,matrix_A[3722],matrix_B[122],mul_res1[3722]);
multi_7x28 multi_7x28_mod_3723(clk,rst,matrix_A[3723],matrix_B[123],mul_res1[3723]);
multi_7x28 multi_7x28_mod_3724(clk,rst,matrix_A[3724],matrix_B[124],mul_res1[3724]);
multi_7x28 multi_7x28_mod_3725(clk,rst,matrix_A[3725],matrix_B[125],mul_res1[3725]);
multi_7x28 multi_7x28_mod_3726(clk,rst,matrix_A[3726],matrix_B[126],mul_res1[3726]);
multi_7x28 multi_7x28_mod_3727(clk,rst,matrix_A[3727],matrix_B[127],mul_res1[3727]);
multi_7x28 multi_7x28_mod_3728(clk,rst,matrix_A[3728],matrix_B[128],mul_res1[3728]);
multi_7x28 multi_7x28_mod_3729(clk,rst,matrix_A[3729],matrix_B[129],mul_res1[3729]);
multi_7x28 multi_7x28_mod_3730(clk,rst,matrix_A[3730],matrix_B[130],mul_res1[3730]);
multi_7x28 multi_7x28_mod_3731(clk,rst,matrix_A[3731],matrix_B[131],mul_res1[3731]);
multi_7x28 multi_7x28_mod_3732(clk,rst,matrix_A[3732],matrix_B[132],mul_res1[3732]);
multi_7x28 multi_7x28_mod_3733(clk,rst,matrix_A[3733],matrix_B[133],mul_res1[3733]);
multi_7x28 multi_7x28_mod_3734(clk,rst,matrix_A[3734],matrix_B[134],mul_res1[3734]);
multi_7x28 multi_7x28_mod_3735(clk,rst,matrix_A[3735],matrix_B[135],mul_res1[3735]);
multi_7x28 multi_7x28_mod_3736(clk,rst,matrix_A[3736],matrix_B[136],mul_res1[3736]);
multi_7x28 multi_7x28_mod_3737(clk,rst,matrix_A[3737],matrix_B[137],mul_res1[3737]);
multi_7x28 multi_7x28_mod_3738(clk,rst,matrix_A[3738],matrix_B[138],mul_res1[3738]);
multi_7x28 multi_7x28_mod_3739(clk,rst,matrix_A[3739],matrix_B[139],mul_res1[3739]);
multi_7x28 multi_7x28_mod_3740(clk,rst,matrix_A[3740],matrix_B[140],mul_res1[3740]);
multi_7x28 multi_7x28_mod_3741(clk,rst,matrix_A[3741],matrix_B[141],mul_res1[3741]);
multi_7x28 multi_7x28_mod_3742(clk,rst,matrix_A[3742],matrix_B[142],mul_res1[3742]);
multi_7x28 multi_7x28_mod_3743(clk,rst,matrix_A[3743],matrix_B[143],mul_res1[3743]);
multi_7x28 multi_7x28_mod_3744(clk,rst,matrix_A[3744],matrix_B[144],mul_res1[3744]);
multi_7x28 multi_7x28_mod_3745(clk,rst,matrix_A[3745],matrix_B[145],mul_res1[3745]);
multi_7x28 multi_7x28_mod_3746(clk,rst,matrix_A[3746],matrix_B[146],mul_res1[3746]);
multi_7x28 multi_7x28_mod_3747(clk,rst,matrix_A[3747],matrix_B[147],mul_res1[3747]);
multi_7x28 multi_7x28_mod_3748(clk,rst,matrix_A[3748],matrix_B[148],mul_res1[3748]);
multi_7x28 multi_7x28_mod_3749(clk,rst,matrix_A[3749],matrix_B[149],mul_res1[3749]);
multi_7x28 multi_7x28_mod_3750(clk,rst,matrix_A[3750],matrix_B[150],mul_res1[3750]);
multi_7x28 multi_7x28_mod_3751(clk,rst,matrix_A[3751],matrix_B[151],mul_res1[3751]);
multi_7x28 multi_7x28_mod_3752(clk,rst,matrix_A[3752],matrix_B[152],mul_res1[3752]);
multi_7x28 multi_7x28_mod_3753(clk,rst,matrix_A[3753],matrix_B[153],mul_res1[3753]);
multi_7x28 multi_7x28_mod_3754(clk,rst,matrix_A[3754],matrix_B[154],mul_res1[3754]);
multi_7x28 multi_7x28_mod_3755(clk,rst,matrix_A[3755],matrix_B[155],mul_res1[3755]);
multi_7x28 multi_7x28_mod_3756(clk,rst,matrix_A[3756],matrix_B[156],mul_res1[3756]);
multi_7x28 multi_7x28_mod_3757(clk,rst,matrix_A[3757],matrix_B[157],mul_res1[3757]);
multi_7x28 multi_7x28_mod_3758(clk,rst,matrix_A[3758],matrix_B[158],mul_res1[3758]);
multi_7x28 multi_7x28_mod_3759(clk,rst,matrix_A[3759],matrix_B[159],mul_res1[3759]);
multi_7x28 multi_7x28_mod_3760(clk,rst,matrix_A[3760],matrix_B[160],mul_res1[3760]);
multi_7x28 multi_7x28_mod_3761(clk,rst,matrix_A[3761],matrix_B[161],mul_res1[3761]);
multi_7x28 multi_7x28_mod_3762(clk,rst,matrix_A[3762],matrix_B[162],mul_res1[3762]);
multi_7x28 multi_7x28_mod_3763(clk,rst,matrix_A[3763],matrix_B[163],mul_res1[3763]);
multi_7x28 multi_7x28_mod_3764(clk,rst,matrix_A[3764],matrix_B[164],mul_res1[3764]);
multi_7x28 multi_7x28_mod_3765(clk,rst,matrix_A[3765],matrix_B[165],mul_res1[3765]);
multi_7x28 multi_7x28_mod_3766(clk,rst,matrix_A[3766],matrix_B[166],mul_res1[3766]);
multi_7x28 multi_7x28_mod_3767(clk,rst,matrix_A[3767],matrix_B[167],mul_res1[3767]);
multi_7x28 multi_7x28_mod_3768(clk,rst,matrix_A[3768],matrix_B[168],mul_res1[3768]);
multi_7x28 multi_7x28_mod_3769(clk,rst,matrix_A[3769],matrix_B[169],mul_res1[3769]);
multi_7x28 multi_7x28_mod_3770(clk,rst,matrix_A[3770],matrix_B[170],mul_res1[3770]);
multi_7x28 multi_7x28_mod_3771(clk,rst,matrix_A[3771],matrix_B[171],mul_res1[3771]);
multi_7x28 multi_7x28_mod_3772(clk,rst,matrix_A[3772],matrix_B[172],mul_res1[3772]);
multi_7x28 multi_7x28_mod_3773(clk,rst,matrix_A[3773],matrix_B[173],mul_res1[3773]);
multi_7x28 multi_7x28_mod_3774(clk,rst,matrix_A[3774],matrix_B[174],mul_res1[3774]);
multi_7x28 multi_7x28_mod_3775(clk,rst,matrix_A[3775],matrix_B[175],mul_res1[3775]);
multi_7x28 multi_7x28_mod_3776(clk,rst,matrix_A[3776],matrix_B[176],mul_res1[3776]);
multi_7x28 multi_7x28_mod_3777(clk,rst,matrix_A[3777],matrix_B[177],mul_res1[3777]);
multi_7x28 multi_7x28_mod_3778(clk,rst,matrix_A[3778],matrix_B[178],mul_res1[3778]);
multi_7x28 multi_7x28_mod_3779(clk,rst,matrix_A[3779],matrix_B[179],mul_res1[3779]);
multi_7x28 multi_7x28_mod_3780(clk,rst,matrix_A[3780],matrix_B[180],mul_res1[3780]);
multi_7x28 multi_7x28_mod_3781(clk,rst,matrix_A[3781],matrix_B[181],mul_res1[3781]);
multi_7x28 multi_7x28_mod_3782(clk,rst,matrix_A[3782],matrix_B[182],mul_res1[3782]);
multi_7x28 multi_7x28_mod_3783(clk,rst,matrix_A[3783],matrix_B[183],mul_res1[3783]);
multi_7x28 multi_7x28_mod_3784(clk,rst,matrix_A[3784],matrix_B[184],mul_res1[3784]);
multi_7x28 multi_7x28_mod_3785(clk,rst,matrix_A[3785],matrix_B[185],mul_res1[3785]);
multi_7x28 multi_7x28_mod_3786(clk,rst,matrix_A[3786],matrix_B[186],mul_res1[3786]);
multi_7x28 multi_7x28_mod_3787(clk,rst,matrix_A[3787],matrix_B[187],mul_res1[3787]);
multi_7x28 multi_7x28_mod_3788(clk,rst,matrix_A[3788],matrix_B[188],mul_res1[3788]);
multi_7x28 multi_7x28_mod_3789(clk,rst,matrix_A[3789],matrix_B[189],mul_res1[3789]);
multi_7x28 multi_7x28_mod_3790(clk,rst,matrix_A[3790],matrix_B[190],mul_res1[3790]);
multi_7x28 multi_7x28_mod_3791(clk,rst,matrix_A[3791],matrix_B[191],mul_res1[3791]);
multi_7x28 multi_7x28_mod_3792(clk,rst,matrix_A[3792],matrix_B[192],mul_res1[3792]);
multi_7x28 multi_7x28_mod_3793(clk,rst,matrix_A[3793],matrix_B[193],mul_res1[3793]);
multi_7x28 multi_7x28_mod_3794(clk,rst,matrix_A[3794],matrix_B[194],mul_res1[3794]);
multi_7x28 multi_7x28_mod_3795(clk,rst,matrix_A[3795],matrix_B[195],mul_res1[3795]);
multi_7x28 multi_7x28_mod_3796(clk,rst,matrix_A[3796],matrix_B[196],mul_res1[3796]);
multi_7x28 multi_7x28_mod_3797(clk,rst,matrix_A[3797],matrix_B[197],mul_res1[3797]);
multi_7x28 multi_7x28_mod_3798(clk,rst,matrix_A[3798],matrix_B[198],mul_res1[3798]);
multi_7x28 multi_7x28_mod_3799(clk,rst,matrix_A[3799],matrix_B[199],mul_res1[3799]);
multi_7x28 multi_7x28_mod_3800(clk,rst,matrix_A[3800],matrix_B[0],mul_res1[3800]);
multi_7x28 multi_7x28_mod_3801(clk,rst,matrix_A[3801],matrix_B[1],mul_res1[3801]);
multi_7x28 multi_7x28_mod_3802(clk,rst,matrix_A[3802],matrix_B[2],mul_res1[3802]);
multi_7x28 multi_7x28_mod_3803(clk,rst,matrix_A[3803],matrix_B[3],mul_res1[3803]);
multi_7x28 multi_7x28_mod_3804(clk,rst,matrix_A[3804],matrix_B[4],mul_res1[3804]);
multi_7x28 multi_7x28_mod_3805(clk,rst,matrix_A[3805],matrix_B[5],mul_res1[3805]);
multi_7x28 multi_7x28_mod_3806(clk,rst,matrix_A[3806],matrix_B[6],mul_res1[3806]);
multi_7x28 multi_7x28_mod_3807(clk,rst,matrix_A[3807],matrix_B[7],mul_res1[3807]);
multi_7x28 multi_7x28_mod_3808(clk,rst,matrix_A[3808],matrix_B[8],mul_res1[3808]);
multi_7x28 multi_7x28_mod_3809(clk,rst,matrix_A[3809],matrix_B[9],mul_res1[3809]);
multi_7x28 multi_7x28_mod_3810(clk,rst,matrix_A[3810],matrix_B[10],mul_res1[3810]);
multi_7x28 multi_7x28_mod_3811(clk,rst,matrix_A[3811],matrix_B[11],mul_res1[3811]);
multi_7x28 multi_7x28_mod_3812(clk,rst,matrix_A[3812],matrix_B[12],mul_res1[3812]);
multi_7x28 multi_7x28_mod_3813(clk,rst,matrix_A[3813],matrix_B[13],mul_res1[3813]);
multi_7x28 multi_7x28_mod_3814(clk,rst,matrix_A[3814],matrix_B[14],mul_res1[3814]);
multi_7x28 multi_7x28_mod_3815(clk,rst,matrix_A[3815],matrix_B[15],mul_res1[3815]);
multi_7x28 multi_7x28_mod_3816(clk,rst,matrix_A[3816],matrix_B[16],mul_res1[3816]);
multi_7x28 multi_7x28_mod_3817(clk,rst,matrix_A[3817],matrix_B[17],mul_res1[3817]);
multi_7x28 multi_7x28_mod_3818(clk,rst,matrix_A[3818],matrix_B[18],mul_res1[3818]);
multi_7x28 multi_7x28_mod_3819(clk,rst,matrix_A[3819],matrix_B[19],mul_res1[3819]);
multi_7x28 multi_7x28_mod_3820(clk,rst,matrix_A[3820],matrix_B[20],mul_res1[3820]);
multi_7x28 multi_7x28_mod_3821(clk,rst,matrix_A[3821],matrix_B[21],mul_res1[3821]);
multi_7x28 multi_7x28_mod_3822(clk,rst,matrix_A[3822],matrix_B[22],mul_res1[3822]);
multi_7x28 multi_7x28_mod_3823(clk,rst,matrix_A[3823],matrix_B[23],mul_res1[3823]);
multi_7x28 multi_7x28_mod_3824(clk,rst,matrix_A[3824],matrix_B[24],mul_res1[3824]);
multi_7x28 multi_7x28_mod_3825(clk,rst,matrix_A[3825],matrix_B[25],mul_res1[3825]);
multi_7x28 multi_7x28_mod_3826(clk,rst,matrix_A[3826],matrix_B[26],mul_res1[3826]);
multi_7x28 multi_7x28_mod_3827(clk,rst,matrix_A[3827],matrix_B[27],mul_res1[3827]);
multi_7x28 multi_7x28_mod_3828(clk,rst,matrix_A[3828],matrix_B[28],mul_res1[3828]);
multi_7x28 multi_7x28_mod_3829(clk,rst,matrix_A[3829],matrix_B[29],mul_res1[3829]);
multi_7x28 multi_7x28_mod_3830(clk,rst,matrix_A[3830],matrix_B[30],mul_res1[3830]);
multi_7x28 multi_7x28_mod_3831(clk,rst,matrix_A[3831],matrix_B[31],mul_res1[3831]);
multi_7x28 multi_7x28_mod_3832(clk,rst,matrix_A[3832],matrix_B[32],mul_res1[3832]);
multi_7x28 multi_7x28_mod_3833(clk,rst,matrix_A[3833],matrix_B[33],mul_res1[3833]);
multi_7x28 multi_7x28_mod_3834(clk,rst,matrix_A[3834],matrix_B[34],mul_res1[3834]);
multi_7x28 multi_7x28_mod_3835(clk,rst,matrix_A[3835],matrix_B[35],mul_res1[3835]);
multi_7x28 multi_7x28_mod_3836(clk,rst,matrix_A[3836],matrix_B[36],mul_res1[3836]);
multi_7x28 multi_7x28_mod_3837(clk,rst,matrix_A[3837],matrix_B[37],mul_res1[3837]);
multi_7x28 multi_7x28_mod_3838(clk,rst,matrix_A[3838],matrix_B[38],mul_res1[3838]);
multi_7x28 multi_7x28_mod_3839(clk,rst,matrix_A[3839],matrix_B[39],mul_res1[3839]);
multi_7x28 multi_7x28_mod_3840(clk,rst,matrix_A[3840],matrix_B[40],mul_res1[3840]);
multi_7x28 multi_7x28_mod_3841(clk,rst,matrix_A[3841],matrix_B[41],mul_res1[3841]);
multi_7x28 multi_7x28_mod_3842(clk,rst,matrix_A[3842],matrix_B[42],mul_res1[3842]);
multi_7x28 multi_7x28_mod_3843(clk,rst,matrix_A[3843],matrix_B[43],mul_res1[3843]);
multi_7x28 multi_7x28_mod_3844(clk,rst,matrix_A[3844],matrix_B[44],mul_res1[3844]);
multi_7x28 multi_7x28_mod_3845(clk,rst,matrix_A[3845],matrix_B[45],mul_res1[3845]);
multi_7x28 multi_7x28_mod_3846(clk,rst,matrix_A[3846],matrix_B[46],mul_res1[3846]);
multi_7x28 multi_7x28_mod_3847(clk,rst,matrix_A[3847],matrix_B[47],mul_res1[3847]);
multi_7x28 multi_7x28_mod_3848(clk,rst,matrix_A[3848],matrix_B[48],mul_res1[3848]);
multi_7x28 multi_7x28_mod_3849(clk,rst,matrix_A[3849],matrix_B[49],mul_res1[3849]);
multi_7x28 multi_7x28_mod_3850(clk,rst,matrix_A[3850],matrix_B[50],mul_res1[3850]);
multi_7x28 multi_7x28_mod_3851(clk,rst,matrix_A[3851],matrix_B[51],mul_res1[3851]);
multi_7x28 multi_7x28_mod_3852(clk,rst,matrix_A[3852],matrix_B[52],mul_res1[3852]);
multi_7x28 multi_7x28_mod_3853(clk,rst,matrix_A[3853],matrix_B[53],mul_res1[3853]);
multi_7x28 multi_7x28_mod_3854(clk,rst,matrix_A[3854],matrix_B[54],mul_res1[3854]);
multi_7x28 multi_7x28_mod_3855(clk,rst,matrix_A[3855],matrix_B[55],mul_res1[3855]);
multi_7x28 multi_7x28_mod_3856(clk,rst,matrix_A[3856],matrix_B[56],mul_res1[3856]);
multi_7x28 multi_7x28_mod_3857(clk,rst,matrix_A[3857],matrix_B[57],mul_res1[3857]);
multi_7x28 multi_7x28_mod_3858(clk,rst,matrix_A[3858],matrix_B[58],mul_res1[3858]);
multi_7x28 multi_7x28_mod_3859(clk,rst,matrix_A[3859],matrix_B[59],mul_res1[3859]);
multi_7x28 multi_7x28_mod_3860(clk,rst,matrix_A[3860],matrix_B[60],mul_res1[3860]);
multi_7x28 multi_7x28_mod_3861(clk,rst,matrix_A[3861],matrix_B[61],mul_res1[3861]);
multi_7x28 multi_7x28_mod_3862(clk,rst,matrix_A[3862],matrix_B[62],mul_res1[3862]);
multi_7x28 multi_7x28_mod_3863(clk,rst,matrix_A[3863],matrix_B[63],mul_res1[3863]);
multi_7x28 multi_7x28_mod_3864(clk,rst,matrix_A[3864],matrix_B[64],mul_res1[3864]);
multi_7x28 multi_7x28_mod_3865(clk,rst,matrix_A[3865],matrix_B[65],mul_res1[3865]);
multi_7x28 multi_7x28_mod_3866(clk,rst,matrix_A[3866],matrix_B[66],mul_res1[3866]);
multi_7x28 multi_7x28_mod_3867(clk,rst,matrix_A[3867],matrix_B[67],mul_res1[3867]);
multi_7x28 multi_7x28_mod_3868(clk,rst,matrix_A[3868],matrix_B[68],mul_res1[3868]);
multi_7x28 multi_7x28_mod_3869(clk,rst,matrix_A[3869],matrix_B[69],mul_res1[3869]);
multi_7x28 multi_7x28_mod_3870(clk,rst,matrix_A[3870],matrix_B[70],mul_res1[3870]);
multi_7x28 multi_7x28_mod_3871(clk,rst,matrix_A[3871],matrix_B[71],mul_res1[3871]);
multi_7x28 multi_7x28_mod_3872(clk,rst,matrix_A[3872],matrix_B[72],mul_res1[3872]);
multi_7x28 multi_7x28_mod_3873(clk,rst,matrix_A[3873],matrix_B[73],mul_res1[3873]);
multi_7x28 multi_7x28_mod_3874(clk,rst,matrix_A[3874],matrix_B[74],mul_res1[3874]);
multi_7x28 multi_7x28_mod_3875(clk,rst,matrix_A[3875],matrix_B[75],mul_res1[3875]);
multi_7x28 multi_7x28_mod_3876(clk,rst,matrix_A[3876],matrix_B[76],mul_res1[3876]);
multi_7x28 multi_7x28_mod_3877(clk,rst,matrix_A[3877],matrix_B[77],mul_res1[3877]);
multi_7x28 multi_7x28_mod_3878(clk,rst,matrix_A[3878],matrix_B[78],mul_res1[3878]);
multi_7x28 multi_7x28_mod_3879(clk,rst,matrix_A[3879],matrix_B[79],mul_res1[3879]);
multi_7x28 multi_7x28_mod_3880(clk,rst,matrix_A[3880],matrix_B[80],mul_res1[3880]);
multi_7x28 multi_7x28_mod_3881(clk,rst,matrix_A[3881],matrix_B[81],mul_res1[3881]);
multi_7x28 multi_7x28_mod_3882(clk,rst,matrix_A[3882],matrix_B[82],mul_res1[3882]);
multi_7x28 multi_7x28_mod_3883(clk,rst,matrix_A[3883],matrix_B[83],mul_res1[3883]);
multi_7x28 multi_7x28_mod_3884(clk,rst,matrix_A[3884],matrix_B[84],mul_res1[3884]);
multi_7x28 multi_7x28_mod_3885(clk,rst,matrix_A[3885],matrix_B[85],mul_res1[3885]);
multi_7x28 multi_7x28_mod_3886(clk,rst,matrix_A[3886],matrix_B[86],mul_res1[3886]);
multi_7x28 multi_7x28_mod_3887(clk,rst,matrix_A[3887],matrix_B[87],mul_res1[3887]);
multi_7x28 multi_7x28_mod_3888(clk,rst,matrix_A[3888],matrix_B[88],mul_res1[3888]);
multi_7x28 multi_7x28_mod_3889(clk,rst,matrix_A[3889],matrix_B[89],mul_res1[3889]);
multi_7x28 multi_7x28_mod_3890(clk,rst,matrix_A[3890],matrix_B[90],mul_res1[3890]);
multi_7x28 multi_7x28_mod_3891(clk,rst,matrix_A[3891],matrix_B[91],mul_res1[3891]);
multi_7x28 multi_7x28_mod_3892(clk,rst,matrix_A[3892],matrix_B[92],mul_res1[3892]);
multi_7x28 multi_7x28_mod_3893(clk,rst,matrix_A[3893],matrix_B[93],mul_res1[3893]);
multi_7x28 multi_7x28_mod_3894(clk,rst,matrix_A[3894],matrix_B[94],mul_res1[3894]);
multi_7x28 multi_7x28_mod_3895(clk,rst,matrix_A[3895],matrix_B[95],mul_res1[3895]);
multi_7x28 multi_7x28_mod_3896(clk,rst,matrix_A[3896],matrix_B[96],mul_res1[3896]);
multi_7x28 multi_7x28_mod_3897(clk,rst,matrix_A[3897],matrix_B[97],mul_res1[3897]);
multi_7x28 multi_7x28_mod_3898(clk,rst,matrix_A[3898],matrix_B[98],mul_res1[3898]);
multi_7x28 multi_7x28_mod_3899(clk,rst,matrix_A[3899],matrix_B[99],mul_res1[3899]);
multi_7x28 multi_7x28_mod_3900(clk,rst,matrix_A[3900],matrix_B[100],mul_res1[3900]);
multi_7x28 multi_7x28_mod_3901(clk,rst,matrix_A[3901],matrix_B[101],mul_res1[3901]);
multi_7x28 multi_7x28_mod_3902(clk,rst,matrix_A[3902],matrix_B[102],mul_res1[3902]);
multi_7x28 multi_7x28_mod_3903(clk,rst,matrix_A[3903],matrix_B[103],mul_res1[3903]);
multi_7x28 multi_7x28_mod_3904(clk,rst,matrix_A[3904],matrix_B[104],mul_res1[3904]);
multi_7x28 multi_7x28_mod_3905(clk,rst,matrix_A[3905],matrix_B[105],mul_res1[3905]);
multi_7x28 multi_7x28_mod_3906(clk,rst,matrix_A[3906],matrix_B[106],mul_res1[3906]);
multi_7x28 multi_7x28_mod_3907(clk,rst,matrix_A[3907],matrix_B[107],mul_res1[3907]);
multi_7x28 multi_7x28_mod_3908(clk,rst,matrix_A[3908],matrix_B[108],mul_res1[3908]);
multi_7x28 multi_7x28_mod_3909(clk,rst,matrix_A[3909],matrix_B[109],mul_res1[3909]);
multi_7x28 multi_7x28_mod_3910(clk,rst,matrix_A[3910],matrix_B[110],mul_res1[3910]);
multi_7x28 multi_7x28_mod_3911(clk,rst,matrix_A[3911],matrix_B[111],mul_res1[3911]);
multi_7x28 multi_7x28_mod_3912(clk,rst,matrix_A[3912],matrix_B[112],mul_res1[3912]);
multi_7x28 multi_7x28_mod_3913(clk,rst,matrix_A[3913],matrix_B[113],mul_res1[3913]);
multi_7x28 multi_7x28_mod_3914(clk,rst,matrix_A[3914],matrix_B[114],mul_res1[3914]);
multi_7x28 multi_7x28_mod_3915(clk,rst,matrix_A[3915],matrix_B[115],mul_res1[3915]);
multi_7x28 multi_7x28_mod_3916(clk,rst,matrix_A[3916],matrix_B[116],mul_res1[3916]);
multi_7x28 multi_7x28_mod_3917(clk,rst,matrix_A[3917],matrix_B[117],mul_res1[3917]);
multi_7x28 multi_7x28_mod_3918(clk,rst,matrix_A[3918],matrix_B[118],mul_res1[3918]);
multi_7x28 multi_7x28_mod_3919(clk,rst,matrix_A[3919],matrix_B[119],mul_res1[3919]);
multi_7x28 multi_7x28_mod_3920(clk,rst,matrix_A[3920],matrix_B[120],mul_res1[3920]);
multi_7x28 multi_7x28_mod_3921(clk,rst,matrix_A[3921],matrix_B[121],mul_res1[3921]);
multi_7x28 multi_7x28_mod_3922(clk,rst,matrix_A[3922],matrix_B[122],mul_res1[3922]);
multi_7x28 multi_7x28_mod_3923(clk,rst,matrix_A[3923],matrix_B[123],mul_res1[3923]);
multi_7x28 multi_7x28_mod_3924(clk,rst,matrix_A[3924],matrix_B[124],mul_res1[3924]);
multi_7x28 multi_7x28_mod_3925(clk,rst,matrix_A[3925],matrix_B[125],mul_res1[3925]);
multi_7x28 multi_7x28_mod_3926(clk,rst,matrix_A[3926],matrix_B[126],mul_res1[3926]);
multi_7x28 multi_7x28_mod_3927(clk,rst,matrix_A[3927],matrix_B[127],mul_res1[3927]);
multi_7x28 multi_7x28_mod_3928(clk,rst,matrix_A[3928],matrix_B[128],mul_res1[3928]);
multi_7x28 multi_7x28_mod_3929(clk,rst,matrix_A[3929],matrix_B[129],mul_res1[3929]);
multi_7x28 multi_7x28_mod_3930(clk,rst,matrix_A[3930],matrix_B[130],mul_res1[3930]);
multi_7x28 multi_7x28_mod_3931(clk,rst,matrix_A[3931],matrix_B[131],mul_res1[3931]);
multi_7x28 multi_7x28_mod_3932(clk,rst,matrix_A[3932],matrix_B[132],mul_res1[3932]);
multi_7x28 multi_7x28_mod_3933(clk,rst,matrix_A[3933],matrix_B[133],mul_res1[3933]);
multi_7x28 multi_7x28_mod_3934(clk,rst,matrix_A[3934],matrix_B[134],mul_res1[3934]);
multi_7x28 multi_7x28_mod_3935(clk,rst,matrix_A[3935],matrix_B[135],mul_res1[3935]);
multi_7x28 multi_7x28_mod_3936(clk,rst,matrix_A[3936],matrix_B[136],mul_res1[3936]);
multi_7x28 multi_7x28_mod_3937(clk,rst,matrix_A[3937],matrix_B[137],mul_res1[3937]);
multi_7x28 multi_7x28_mod_3938(clk,rst,matrix_A[3938],matrix_B[138],mul_res1[3938]);
multi_7x28 multi_7x28_mod_3939(clk,rst,matrix_A[3939],matrix_B[139],mul_res1[3939]);
multi_7x28 multi_7x28_mod_3940(clk,rst,matrix_A[3940],matrix_B[140],mul_res1[3940]);
multi_7x28 multi_7x28_mod_3941(clk,rst,matrix_A[3941],matrix_B[141],mul_res1[3941]);
multi_7x28 multi_7x28_mod_3942(clk,rst,matrix_A[3942],matrix_B[142],mul_res1[3942]);
multi_7x28 multi_7x28_mod_3943(clk,rst,matrix_A[3943],matrix_B[143],mul_res1[3943]);
multi_7x28 multi_7x28_mod_3944(clk,rst,matrix_A[3944],matrix_B[144],mul_res1[3944]);
multi_7x28 multi_7x28_mod_3945(clk,rst,matrix_A[3945],matrix_B[145],mul_res1[3945]);
multi_7x28 multi_7x28_mod_3946(clk,rst,matrix_A[3946],matrix_B[146],mul_res1[3946]);
multi_7x28 multi_7x28_mod_3947(clk,rst,matrix_A[3947],matrix_B[147],mul_res1[3947]);
multi_7x28 multi_7x28_mod_3948(clk,rst,matrix_A[3948],matrix_B[148],mul_res1[3948]);
multi_7x28 multi_7x28_mod_3949(clk,rst,matrix_A[3949],matrix_B[149],mul_res1[3949]);
multi_7x28 multi_7x28_mod_3950(clk,rst,matrix_A[3950],matrix_B[150],mul_res1[3950]);
multi_7x28 multi_7x28_mod_3951(clk,rst,matrix_A[3951],matrix_B[151],mul_res1[3951]);
multi_7x28 multi_7x28_mod_3952(clk,rst,matrix_A[3952],matrix_B[152],mul_res1[3952]);
multi_7x28 multi_7x28_mod_3953(clk,rst,matrix_A[3953],matrix_B[153],mul_res1[3953]);
multi_7x28 multi_7x28_mod_3954(clk,rst,matrix_A[3954],matrix_B[154],mul_res1[3954]);
multi_7x28 multi_7x28_mod_3955(clk,rst,matrix_A[3955],matrix_B[155],mul_res1[3955]);
multi_7x28 multi_7x28_mod_3956(clk,rst,matrix_A[3956],matrix_B[156],mul_res1[3956]);
multi_7x28 multi_7x28_mod_3957(clk,rst,matrix_A[3957],matrix_B[157],mul_res1[3957]);
multi_7x28 multi_7x28_mod_3958(clk,rst,matrix_A[3958],matrix_B[158],mul_res1[3958]);
multi_7x28 multi_7x28_mod_3959(clk,rst,matrix_A[3959],matrix_B[159],mul_res1[3959]);
multi_7x28 multi_7x28_mod_3960(clk,rst,matrix_A[3960],matrix_B[160],mul_res1[3960]);
multi_7x28 multi_7x28_mod_3961(clk,rst,matrix_A[3961],matrix_B[161],mul_res1[3961]);
multi_7x28 multi_7x28_mod_3962(clk,rst,matrix_A[3962],matrix_B[162],mul_res1[3962]);
multi_7x28 multi_7x28_mod_3963(clk,rst,matrix_A[3963],matrix_B[163],mul_res1[3963]);
multi_7x28 multi_7x28_mod_3964(clk,rst,matrix_A[3964],matrix_B[164],mul_res1[3964]);
multi_7x28 multi_7x28_mod_3965(clk,rst,matrix_A[3965],matrix_B[165],mul_res1[3965]);
multi_7x28 multi_7x28_mod_3966(clk,rst,matrix_A[3966],matrix_B[166],mul_res1[3966]);
multi_7x28 multi_7x28_mod_3967(clk,rst,matrix_A[3967],matrix_B[167],mul_res1[3967]);
multi_7x28 multi_7x28_mod_3968(clk,rst,matrix_A[3968],matrix_B[168],mul_res1[3968]);
multi_7x28 multi_7x28_mod_3969(clk,rst,matrix_A[3969],matrix_B[169],mul_res1[3969]);
multi_7x28 multi_7x28_mod_3970(clk,rst,matrix_A[3970],matrix_B[170],mul_res1[3970]);
multi_7x28 multi_7x28_mod_3971(clk,rst,matrix_A[3971],matrix_B[171],mul_res1[3971]);
multi_7x28 multi_7x28_mod_3972(clk,rst,matrix_A[3972],matrix_B[172],mul_res1[3972]);
multi_7x28 multi_7x28_mod_3973(clk,rst,matrix_A[3973],matrix_B[173],mul_res1[3973]);
multi_7x28 multi_7x28_mod_3974(clk,rst,matrix_A[3974],matrix_B[174],mul_res1[3974]);
multi_7x28 multi_7x28_mod_3975(clk,rst,matrix_A[3975],matrix_B[175],mul_res1[3975]);
multi_7x28 multi_7x28_mod_3976(clk,rst,matrix_A[3976],matrix_B[176],mul_res1[3976]);
multi_7x28 multi_7x28_mod_3977(clk,rst,matrix_A[3977],matrix_B[177],mul_res1[3977]);
multi_7x28 multi_7x28_mod_3978(clk,rst,matrix_A[3978],matrix_B[178],mul_res1[3978]);
multi_7x28 multi_7x28_mod_3979(clk,rst,matrix_A[3979],matrix_B[179],mul_res1[3979]);
multi_7x28 multi_7x28_mod_3980(clk,rst,matrix_A[3980],matrix_B[180],mul_res1[3980]);
multi_7x28 multi_7x28_mod_3981(clk,rst,matrix_A[3981],matrix_B[181],mul_res1[3981]);
multi_7x28 multi_7x28_mod_3982(clk,rst,matrix_A[3982],matrix_B[182],mul_res1[3982]);
multi_7x28 multi_7x28_mod_3983(clk,rst,matrix_A[3983],matrix_B[183],mul_res1[3983]);
multi_7x28 multi_7x28_mod_3984(clk,rst,matrix_A[3984],matrix_B[184],mul_res1[3984]);
multi_7x28 multi_7x28_mod_3985(clk,rst,matrix_A[3985],matrix_B[185],mul_res1[3985]);
multi_7x28 multi_7x28_mod_3986(clk,rst,matrix_A[3986],matrix_B[186],mul_res1[3986]);
multi_7x28 multi_7x28_mod_3987(clk,rst,matrix_A[3987],matrix_B[187],mul_res1[3987]);
multi_7x28 multi_7x28_mod_3988(clk,rst,matrix_A[3988],matrix_B[188],mul_res1[3988]);
multi_7x28 multi_7x28_mod_3989(clk,rst,matrix_A[3989],matrix_B[189],mul_res1[3989]);
multi_7x28 multi_7x28_mod_3990(clk,rst,matrix_A[3990],matrix_B[190],mul_res1[3990]);
multi_7x28 multi_7x28_mod_3991(clk,rst,matrix_A[3991],matrix_B[191],mul_res1[3991]);
multi_7x28 multi_7x28_mod_3992(clk,rst,matrix_A[3992],matrix_B[192],mul_res1[3992]);
multi_7x28 multi_7x28_mod_3993(clk,rst,matrix_A[3993],matrix_B[193],mul_res1[3993]);
multi_7x28 multi_7x28_mod_3994(clk,rst,matrix_A[3994],matrix_B[194],mul_res1[3994]);
multi_7x28 multi_7x28_mod_3995(clk,rst,matrix_A[3995],matrix_B[195],mul_res1[3995]);
multi_7x28 multi_7x28_mod_3996(clk,rst,matrix_A[3996],matrix_B[196],mul_res1[3996]);
multi_7x28 multi_7x28_mod_3997(clk,rst,matrix_A[3997],matrix_B[197],mul_res1[3997]);
multi_7x28 multi_7x28_mod_3998(clk,rst,matrix_A[3998],matrix_B[198],mul_res1[3998]);
multi_7x28 multi_7x28_mod_3999(clk,rst,matrix_A[3999],matrix_B[199],mul_res1[3999]);
multi_7x28 multi_7x28_mod_4000(clk,rst,matrix_A[4000],matrix_B[0],mul_res1[4000]);
multi_7x28 multi_7x28_mod_4001(clk,rst,matrix_A[4001],matrix_B[1],mul_res1[4001]);
multi_7x28 multi_7x28_mod_4002(clk,rst,matrix_A[4002],matrix_B[2],mul_res1[4002]);
multi_7x28 multi_7x28_mod_4003(clk,rst,matrix_A[4003],matrix_B[3],mul_res1[4003]);
multi_7x28 multi_7x28_mod_4004(clk,rst,matrix_A[4004],matrix_B[4],mul_res1[4004]);
multi_7x28 multi_7x28_mod_4005(clk,rst,matrix_A[4005],matrix_B[5],mul_res1[4005]);
multi_7x28 multi_7x28_mod_4006(clk,rst,matrix_A[4006],matrix_B[6],mul_res1[4006]);
multi_7x28 multi_7x28_mod_4007(clk,rst,matrix_A[4007],matrix_B[7],mul_res1[4007]);
multi_7x28 multi_7x28_mod_4008(clk,rst,matrix_A[4008],matrix_B[8],mul_res1[4008]);
multi_7x28 multi_7x28_mod_4009(clk,rst,matrix_A[4009],matrix_B[9],mul_res1[4009]);
multi_7x28 multi_7x28_mod_4010(clk,rst,matrix_A[4010],matrix_B[10],mul_res1[4010]);
multi_7x28 multi_7x28_mod_4011(clk,rst,matrix_A[4011],matrix_B[11],mul_res1[4011]);
multi_7x28 multi_7x28_mod_4012(clk,rst,matrix_A[4012],matrix_B[12],mul_res1[4012]);
multi_7x28 multi_7x28_mod_4013(clk,rst,matrix_A[4013],matrix_B[13],mul_res1[4013]);
multi_7x28 multi_7x28_mod_4014(clk,rst,matrix_A[4014],matrix_B[14],mul_res1[4014]);
multi_7x28 multi_7x28_mod_4015(clk,rst,matrix_A[4015],matrix_B[15],mul_res1[4015]);
multi_7x28 multi_7x28_mod_4016(clk,rst,matrix_A[4016],matrix_B[16],mul_res1[4016]);
multi_7x28 multi_7x28_mod_4017(clk,rst,matrix_A[4017],matrix_B[17],mul_res1[4017]);
multi_7x28 multi_7x28_mod_4018(clk,rst,matrix_A[4018],matrix_B[18],mul_res1[4018]);
multi_7x28 multi_7x28_mod_4019(clk,rst,matrix_A[4019],matrix_B[19],mul_res1[4019]);
multi_7x28 multi_7x28_mod_4020(clk,rst,matrix_A[4020],matrix_B[20],mul_res1[4020]);
multi_7x28 multi_7x28_mod_4021(clk,rst,matrix_A[4021],matrix_B[21],mul_res1[4021]);
multi_7x28 multi_7x28_mod_4022(clk,rst,matrix_A[4022],matrix_B[22],mul_res1[4022]);
multi_7x28 multi_7x28_mod_4023(clk,rst,matrix_A[4023],matrix_B[23],mul_res1[4023]);
multi_7x28 multi_7x28_mod_4024(clk,rst,matrix_A[4024],matrix_B[24],mul_res1[4024]);
multi_7x28 multi_7x28_mod_4025(clk,rst,matrix_A[4025],matrix_B[25],mul_res1[4025]);
multi_7x28 multi_7x28_mod_4026(clk,rst,matrix_A[4026],matrix_B[26],mul_res1[4026]);
multi_7x28 multi_7x28_mod_4027(clk,rst,matrix_A[4027],matrix_B[27],mul_res1[4027]);
multi_7x28 multi_7x28_mod_4028(clk,rst,matrix_A[4028],matrix_B[28],mul_res1[4028]);
multi_7x28 multi_7x28_mod_4029(clk,rst,matrix_A[4029],matrix_B[29],mul_res1[4029]);
multi_7x28 multi_7x28_mod_4030(clk,rst,matrix_A[4030],matrix_B[30],mul_res1[4030]);
multi_7x28 multi_7x28_mod_4031(clk,rst,matrix_A[4031],matrix_B[31],mul_res1[4031]);
multi_7x28 multi_7x28_mod_4032(clk,rst,matrix_A[4032],matrix_B[32],mul_res1[4032]);
multi_7x28 multi_7x28_mod_4033(clk,rst,matrix_A[4033],matrix_B[33],mul_res1[4033]);
multi_7x28 multi_7x28_mod_4034(clk,rst,matrix_A[4034],matrix_B[34],mul_res1[4034]);
multi_7x28 multi_7x28_mod_4035(clk,rst,matrix_A[4035],matrix_B[35],mul_res1[4035]);
multi_7x28 multi_7x28_mod_4036(clk,rst,matrix_A[4036],matrix_B[36],mul_res1[4036]);
multi_7x28 multi_7x28_mod_4037(clk,rst,matrix_A[4037],matrix_B[37],mul_res1[4037]);
multi_7x28 multi_7x28_mod_4038(clk,rst,matrix_A[4038],matrix_B[38],mul_res1[4038]);
multi_7x28 multi_7x28_mod_4039(clk,rst,matrix_A[4039],matrix_B[39],mul_res1[4039]);
multi_7x28 multi_7x28_mod_4040(clk,rst,matrix_A[4040],matrix_B[40],mul_res1[4040]);
multi_7x28 multi_7x28_mod_4041(clk,rst,matrix_A[4041],matrix_B[41],mul_res1[4041]);
multi_7x28 multi_7x28_mod_4042(clk,rst,matrix_A[4042],matrix_B[42],mul_res1[4042]);
multi_7x28 multi_7x28_mod_4043(clk,rst,matrix_A[4043],matrix_B[43],mul_res1[4043]);
multi_7x28 multi_7x28_mod_4044(clk,rst,matrix_A[4044],matrix_B[44],mul_res1[4044]);
multi_7x28 multi_7x28_mod_4045(clk,rst,matrix_A[4045],matrix_B[45],mul_res1[4045]);
multi_7x28 multi_7x28_mod_4046(clk,rst,matrix_A[4046],matrix_B[46],mul_res1[4046]);
multi_7x28 multi_7x28_mod_4047(clk,rst,matrix_A[4047],matrix_B[47],mul_res1[4047]);
multi_7x28 multi_7x28_mod_4048(clk,rst,matrix_A[4048],matrix_B[48],mul_res1[4048]);
multi_7x28 multi_7x28_mod_4049(clk,rst,matrix_A[4049],matrix_B[49],mul_res1[4049]);
multi_7x28 multi_7x28_mod_4050(clk,rst,matrix_A[4050],matrix_B[50],mul_res1[4050]);
multi_7x28 multi_7x28_mod_4051(clk,rst,matrix_A[4051],matrix_B[51],mul_res1[4051]);
multi_7x28 multi_7x28_mod_4052(clk,rst,matrix_A[4052],matrix_B[52],mul_res1[4052]);
multi_7x28 multi_7x28_mod_4053(clk,rst,matrix_A[4053],matrix_B[53],mul_res1[4053]);
multi_7x28 multi_7x28_mod_4054(clk,rst,matrix_A[4054],matrix_B[54],mul_res1[4054]);
multi_7x28 multi_7x28_mod_4055(clk,rst,matrix_A[4055],matrix_B[55],mul_res1[4055]);
multi_7x28 multi_7x28_mod_4056(clk,rst,matrix_A[4056],matrix_B[56],mul_res1[4056]);
multi_7x28 multi_7x28_mod_4057(clk,rst,matrix_A[4057],matrix_B[57],mul_res1[4057]);
multi_7x28 multi_7x28_mod_4058(clk,rst,matrix_A[4058],matrix_B[58],mul_res1[4058]);
multi_7x28 multi_7x28_mod_4059(clk,rst,matrix_A[4059],matrix_B[59],mul_res1[4059]);
multi_7x28 multi_7x28_mod_4060(clk,rst,matrix_A[4060],matrix_B[60],mul_res1[4060]);
multi_7x28 multi_7x28_mod_4061(clk,rst,matrix_A[4061],matrix_B[61],mul_res1[4061]);
multi_7x28 multi_7x28_mod_4062(clk,rst,matrix_A[4062],matrix_B[62],mul_res1[4062]);
multi_7x28 multi_7x28_mod_4063(clk,rst,matrix_A[4063],matrix_B[63],mul_res1[4063]);
multi_7x28 multi_7x28_mod_4064(clk,rst,matrix_A[4064],matrix_B[64],mul_res1[4064]);
multi_7x28 multi_7x28_mod_4065(clk,rst,matrix_A[4065],matrix_B[65],mul_res1[4065]);
multi_7x28 multi_7x28_mod_4066(clk,rst,matrix_A[4066],matrix_B[66],mul_res1[4066]);
multi_7x28 multi_7x28_mod_4067(clk,rst,matrix_A[4067],matrix_B[67],mul_res1[4067]);
multi_7x28 multi_7x28_mod_4068(clk,rst,matrix_A[4068],matrix_B[68],mul_res1[4068]);
multi_7x28 multi_7x28_mod_4069(clk,rst,matrix_A[4069],matrix_B[69],mul_res1[4069]);
multi_7x28 multi_7x28_mod_4070(clk,rst,matrix_A[4070],matrix_B[70],mul_res1[4070]);
multi_7x28 multi_7x28_mod_4071(clk,rst,matrix_A[4071],matrix_B[71],mul_res1[4071]);
multi_7x28 multi_7x28_mod_4072(clk,rst,matrix_A[4072],matrix_B[72],mul_res1[4072]);
multi_7x28 multi_7x28_mod_4073(clk,rst,matrix_A[4073],matrix_B[73],mul_res1[4073]);
multi_7x28 multi_7x28_mod_4074(clk,rst,matrix_A[4074],matrix_B[74],mul_res1[4074]);
multi_7x28 multi_7x28_mod_4075(clk,rst,matrix_A[4075],matrix_B[75],mul_res1[4075]);
multi_7x28 multi_7x28_mod_4076(clk,rst,matrix_A[4076],matrix_B[76],mul_res1[4076]);
multi_7x28 multi_7x28_mod_4077(clk,rst,matrix_A[4077],matrix_B[77],mul_res1[4077]);
multi_7x28 multi_7x28_mod_4078(clk,rst,matrix_A[4078],matrix_B[78],mul_res1[4078]);
multi_7x28 multi_7x28_mod_4079(clk,rst,matrix_A[4079],matrix_B[79],mul_res1[4079]);
multi_7x28 multi_7x28_mod_4080(clk,rst,matrix_A[4080],matrix_B[80],mul_res1[4080]);
multi_7x28 multi_7x28_mod_4081(clk,rst,matrix_A[4081],matrix_B[81],mul_res1[4081]);
multi_7x28 multi_7x28_mod_4082(clk,rst,matrix_A[4082],matrix_B[82],mul_res1[4082]);
multi_7x28 multi_7x28_mod_4083(clk,rst,matrix_A[4083],matrix_B[83],mul_res1[4083]);
multi_7x28 multi_7x28_mod_4084(clk,rst,matrix_A[4084],matrix_B[84],mul_res1[4084]);
multi_7x28 multi_7x28_mod_4085(clk,rst,matrix_A[4085],matrix_B[85],mul_res1[4085]);
multi_7x28 multi_7x28_mod_4086(clk,rst,matrix_A[4086],matrix_B[86],mul_res1[4086]);
multi_7x28 multi_7x28_mod_4087(clk,rst,matrix_A[4087],matrix_B[87],mul_res1[4087]);
multi_7x28 multi_7x28_mod_4088(clk,rst,matrix_A[4088],matrix_B[88],mul_res1[4088]);
multi_7x28 multi_7x28_mod_4089(clk,rst,matrix_A[4089],matrix_B[89],mul_res1[4089]);
multi_7x28 multi_7x28_mod_4090(clk,rst,matrix_A[4090],matrix_B[90],mul_res1[4090]);
multi_7x28 multi_7x28_mod_4091(clk,rst,matrix_A[4091],matrix_B[91],mul_res1[4091]);
multi_7x28 multi_7x28_mod_4092(clk,rst,matrix_A[4092],matrix_B[92],mul_res1[4092]);
multi_7x28 multi_7x28_mod_4093(clk,rst,matrix_A[4093],matrix_B[93],mul_res1[4093]);
multi_7x28 multi_7x28_mod_4094(clk,rst,matrix_A[4094],matrix_B[94],mul_res1[4094]);
multi_7x28 multi_7x28_mod_4095(clk,rst,matrix_A[4095],matrix_B[95],mul_res1[4095]);
multi_7x28 multi_7x28_mod_4096(clk,rst,matrix_A[4096],matrix_B[96],mul_res1[4096]);
multi_7x28 multi_7x28_mod_4097(clk,rst,matrix_A[4097],matrix_B[97],mul_res1[4097]);
multi_7x28 multi_7x28_mod_4098(clk,rst,matrix_A[4098],matrix_B[98],mul_res1[4098]);
multi_7x28 multi_7x28_mod_4099(clk,rst,matrix_A[4099],matrix_B[99],mul_res1[4099]);
multi_7x28 multi_7x28_mod_4100(clk,rst,matrix_A[4100],matrix_B[100],mul_res1[4100]);
multi_7x28 multi_7x28_mod_4101(clk,rst,matrix_A[4101],matrix_B[101],mul_res1[4101]);
multi_7x28 multi_7x28_mod_4102(clk,rst,matrix_A[4102],matrix_B[102],mul_res1[4102]);
multi_7x28 multi_7x28_mod_4103(clk,rst,matrix_A[4103],matrix_B[103],mul_res1[4103]);
multi_7x28 multi_7x28_mod_4104(clk,rst,matrix_A[4104],matrix_B[104],mul_res1[4104]);
multi_7x28 multi_7x28_mod_4105(clk,rst,matrix_A[4105],matrix_B[105],mul_res1[4105]);
multi_7x28 multi_7x28_mod_4106(clk,rst,matrix_A[4106],matrix_B[106],mul_res1[4106]);
multi_7x28 multi_7x28_mod_4107(clk,rst,matrix_A[4107],matrix_B[107],mul_res1[4107]);
multi_7x28 multi_7x28_mod_4108(clk,rst,matrix_A[4108],matrix_B[108],mul_res1[4108]);
multi_7x28 multi_7x28_mod_4109(clk,rst,matrix_A[4109],matrix_B[109],mul_res1[4109]);
multi_7x28 multi_7x28_mod_4110(clk,rst,matrix_A[4110],matrix_B[110],mul_res1[4110]);
multi_7x28 multi_7x28_mod_4111(clk,rst,matrix_A[4111],matrix_B[111],mul_res1[4111]);
multi_7x28 multi_7x28_mod_4112(clk,rst,matrix_A[4112],matrix_B[112],mul_res1[4112]);
multi_7x28 multi_7x28_mod_4113(clk,rst,matrix_A[4113],matrix_B[113],mul_res1[4113]);
multi_7x28 multi_7x28_mod_4114(clk,rst,matrix_A[4114],matrix_B[114],mul_res1[4114]);
multi_7x28 multi_7x28_mod_4115(clk,rst,matrix_A[4115],matrix_B[115],mul_res1[4115]);
multi_7x28 multi_7x28_mod_4116(clk,rst,matrix_A[4116],matrix_B[116],mul_res1[4116]);
multi_7x28 multi_7x28_mod_4117(clk,rst,matrix_A[4117],matrix_B[117],mul_res1[4117]);
multi_7x28 multi_7x28_mod_4118(clk,rst,matrix_A[4118],matrix_B[118],mul_res1[4118]);
multi_7x28 multi_7x28_mod_4119(clk,rst,matrix_A[4119],matrix_B[119],mul_res1[4119]);
multi_7x28 multi_7x28_mod_4120(clk,rst,matrix_A[4120],matrix_B[120],mul_res1[4120]);
multi_7x28 multi_7x28_mod_4121(clk,rst,matrix_A[4121],matrix_B[121],mul_res1[4121]);
multi_7x28 multi_7x28_mod_4122(clk,rst,matrix_A[4122],matrix_B[122],mul_res1[4122]);
multi_7x28 multi_7x28_mod_4123(clk,rst,matrix_A[4123],matrix_B[123],mul_res1[4123]);
multi_7x28 multi_7x28_mod_4124(clk,rst,matrix_A[4124],matrix_B[124],mul_res1[4124]);
multi_7x28 multi_7x28_mod_4125(clk,rst,matrix_A[4125],matrix_B[125],mul_res1[4125]);
multi_7x28 multi_7x28_mod_4126(clk,rst,matrix_A[4126],matrix_B[126],mul_res1[4126]);
multi_7x28 multi_7x28_mod_4127(clk,rst,matrix_A[4127],matrix_B[127],mul_res1[4127]);
multi_7x28 multi_7x28_mod_4128(clk,rst,matrix_A[4128],matrix_B[128],mul_res1[4128]);
multi_7x28 multi_7x28_mod_4129(clk,rst,matrix_A[4129],matrix_B[129],mul_res1[4129]);
multi_7x28 multi_7x28_mod_4130(clk,rst,matrix_A[4130],matrix_B[130],mul_res1[4130]);
multi_7x28 multi_7x28_mod_4131(clk,rst,matrix_A[4131],matrix_B[131],mul_res1[4131]);
multi_7x28 multi_7x28_mod_4132(clk,rst,matrix_A[4132],matrix_B[132],mul_res1[4132]);
multi_7x28 multi_7x28_mod_4133(clk,rst,matrix_A[4133],matrix_B[133],mul_res1[4133]);
multi_7x28 multi_7x28_mod_4134(clk,rst,matrix_A[4134],matrix_B[134],mul_res1[4134]);
multi_7x28 multi_7x28_mod_4135(clk,rst,matrix_A[4135],matrix_B[135],mul_res1[4135]);
multi_7x28 multi_7x28_mod_4136(clk,rst,matrix_A[4136],matrix_B[136],mul_res1[4136]);
multi_7x28 multi_7x28_mod_4137(clk,rst,matrix_A[4137],matrix_B[137],mul_res1[4137]);
multi_7x28 multi_7x28_mod_4138(clk,rst,matrix_A[4138],matrix_B[138],mul_res1[4138]);
multi_7x28 multi_7x28_mod_4139(clk,rst,matrix_A[4139],matrix_B[139],mul_res1[4139]);
multi_7x28 multi_7x28_mod_4140(clk,rst,matrix_A[4140],matrix_B[140],mul_res1[4140]);
multi_7x28 multi_7x28_mod_4141(clk,rst,matrix_A[4141],matrix_B[141],mul_res1[4141]);
multi_7x28 multi_7x28_mod_4142(clk,rst,matrix_A[4142],matrix_B[142],mul_res1[4142]);
multi_7x28 multi_7x28_mod_4143(clk,rst,matrix_A[4143],matrix_B[143],mul_res1[4143]);
multi_7x28 multi_7x28_mod_4144(clk,rst,matrix_A[4144],matrix_B[144],mul_res1[4144]);
multi_7x28 multi_7x28_mod_4145(clk,rst,matrix_A[4145],matrix_B[145],mul_res1[4145]);
multi_7x28 multi_7x28_mod_4146(clk,rst,matrix_A[4146],matrix_B[146],mul_res1[4146]);
multi_7x28 multi_7x28_mod_4147(clk,rst,matrix_A[4147],matrix_B[147],mul_res1[4147]);
multi_7x28 multi_7x28_mod_4148(clk,rst,matrix_A[4148],matrix_B[148],mul_res1[4148]);
multi_7x28 multi_7x28_mod_4149(clk,rst,matrix_A[4149],matrix_B[149],mul_res1[4149]);
multi_7x28 multi_7x28_mod_4150(clk,rst,matrix_A[4150],matrix_B[150],mul_res1[4150]);
multi_7x28 multi_7x28_mod_4151(clk,rst,matrix_A[4151],matrix_B[151],mul_res1[4151]);
multi_7x28 multi_7x28_mod_4152(clk,rst,matrix_A[4152],matrix_B[152],mul_res1[4152]);
multi_7x28 multi_7x28_mod_4153(clk,rst,matrix_A[4153],matrix_B[153],mul_res1[4153]);
multi_7x28 multi_7x28_mod_4154(clk,rst,matrix_A[4154],matrix_B[154],mul_res1[4154]);
multi_7x28 multi_7x28_mod_4155(clk,rst,matrix_A[4155],matrix_B[155],mul_res1[4155]);
multi_7x28 multi_7x28_mod_4156(clk,rst,matrix_A[4156],matrix_B[156],mul_res1[4156]);
multi_7x28 multi_7x28_mod_4157(clk,rst,matrix_A[4157],matrix_B[157],mul_res1[4157]);
multi_7x28 multi_7x28_mod_4158(clk,rst,matrix_A[4158],matrix_B[158],mul_res1[4158]);
multi_7x28 multi_7x28_mod_4159(clk,rst,matrix_A[4159],matrix_B[159],mul_res1[4159]);
multi_7x28 multi_7x28_mod_4160(clk,rst,matrix_A[4160],matrix_B[160],mul_res1[4160]);
multi_7x28 multi_7x28_mod_4161(clk,rst,matrix_A[4161],matrix_B[161],mul_res1[4161]);
multi_7x28 multi_7x28_mod_4162(clk,rst,matrix_A[4162],matrix_B[162],mul_res1[4162]);
multi_7x28 multi_7x28_mod_4163(clk,rst,matrix_A[4163],matrix_B[163],mul_res1[4163]);
multi_7x28 multi_7x28_mod_4164(clk,rst,matrix_A[4164],matrix_B[164],mul_res1[4164]);
multi_7x28 multi_7x28_mod_4165(clk,rst,matrix_A[4165],matrix_B[165],mul_res1[4165]);
multi_7x28 multi_7x28_mod_4166(clk,rst,matrix_A[4166],matrix_B[166],mul_res1[4166]);
multi_7x28 multi_7x28_mod_4167(clk,rst,matrix_A[4167],matrix_B[167],mul_res1[4167]);
multi_7x28 multi_7x28_mod_4168(clk,rst,matrix_A[4168],matrix_B[168],mul_res1[4168]);
multi_7x28 multi_7x28_mod_4169(clk,rst,matrix_A[4169],matrix_B[169],mul_res1[4169]);
multi_7x28 multi_7x28_mod_4170(clk,rst,matrix_A[4170],matrix_B[170],mul_res1[4170]);
multi_7x28 multi_7x28_mod_4171(clk,rst,matrix_A[4171],matrix_B[171],mul_res1[4171]);
multi_7x28 multi_7x28_mod_4172(clk,rst,matrix_A[4172],matrix_B[172],mul_res1[4172]);
multi_7x28 multi_7x28_mod_4173(clk,rst,matrix_A[4173],matrix_B[173],mul_res1[4173]);
multi_7x28 multi_7x28_mod_4174(clk,rst,matrix_A[4174],matrix_B[174],mul_res1[4174]);
multi_7x28 multi_7x28_mod_4175(clk,rst,matrix_A[4175],matrix_B[175],mul_res1[4175]);
multi_7x28 multi_7x28_mod_4176(clk,rst,matrix_A[4176],matrix_B[176],mul_res1[4176]);
multi_7x28 multi_7x28_mod_4177(clk,rst,matrix_A[4177],matrix_B[177],mul_res1[4177]);
multi_7x28 multi_7x28_mod_4178(clk,rst,matrix_A[4178],matrix_B[178],mul_res1[4178]);
multi_7x28 multi_7x28_mod_4179(clk,rst,matrix_A[4179],matrix_B[179],mul_res1[4179]);
multi_7x28 multi_7x28_mod_4180(clk,rst,matrix_A[4180],matrix_B[180],mul_res1[4180]);
multi_7x28 multi_7x28_mod_4181(clk,rst,matrix_A[4181],matrix_B[181],mul_res1[4181]);
multi_7x28 multi_7x28_mod_4182(clk,rst,matrix_A[4182],matrix_B[182],mul_res1[4182]);
multi_7x28 multi_7x28_mod_4183(clk,rst,matrix_A[4183],matrix_B[183],mul_res1[4183]);
multi_7x28 multi_7x28_mod_4184(clk,rst,matrix_A[4184],matrix_B[184],mul_res1[4184]);
multi_7x28 multi_7x28_mod_4185(clk,rst,matrix_A[4185],matrix_B[185],mul_res1[4185]);
multi_7x28 multi_7x28_mod_4186(clk,rst,matrix_A[4186],matrix_B[186],mul_res1[4186]);
multi_7x28 multi_7x28_mod_4187(clk,rst,matrix_A[4187],matrix_B[187],mul_res1[4187]);
multi_7x28 multi_7x28_mod_4188(clk,rst,matrix_A[4188],matrix_B[188],mul_res1[4188]);
multi_7x28 multi_7x28_mod_4189(clk,rst,matrix_A[4189],matrix_B[189],mul_res1[4189]);
multi_7x28 multi_7x28_mod_4190(clk,rst,matrix_A[4190],matrix_B[190],mul_res1[4190]);
multi_7x28 multi_7x28_mod_4191(clk,rst,matrix_A[4191],matrix_B[191],mul_res1[4191]);
multi_7x28 multi_7x28_mod_4192(clk,rst,matrix_A[4192],matrix_B[192],mul_res1[4192]);
multi_7x28 multi_7x28_mod_4193(clk,rst,matrix_A[4193],matrix_B[193],mul_res1[4193]);
multi_7x28 multi_7x28_mod_4194(clk,rst,matrix_A[4194],matrix_B[194],mul_res1[4194]);
multi_7x28 multi_7x28_mod_4195(clk,rst,matrix_A[4195],matrix_B[195],mul_res1[4195]);
multi_7x28 multi_7x28_mod_4196(clk,rst,matrix_A[4196],matrix_B[196],mul_res1[4196]);
multi_7x28 multi_7x28_mod_4197(clk,rst,matrix_A[4197],matrix_B[197],mul_res1[4197]);
multi_7x28 multi_7x28_mod_4198(clk,rst,matrix_A[4198],matrix_B[198],mul_res1[4198]);
multi_7x28 multi_7x28_mod_4199(clk,rst,matrix_A[4199],matrix_B[199],mul_res1[4199]);
multi_7x28 multi_7x28_mod_4200(clk,rst,matrix_A[4200],matrix_B[0],mul_res1[4200]);
multi_7x28 multi_7x28_mod_4201(clk,rst,matrix_A[4201],matrix_B[1],mul_res1[4201]);
multi_7x28 multi_7x28_mod_4202(clk,rst,matrix_A[4202],matrix_B[2],mul_res1[4202]);
multi_7x28 multi_7x28_mod_4203(clk,rst,matrix_A[4203],matrix_B[3],mul_res1[4203]);
multi_7x28 multi_7x28_mod_4204(clk,rst,matrix_A[4204],matrix_B[4],mul_res1[4204]);
multi_7x28 multi_7x28_mod_4205(clk,rst,matrix_A[4205],matrix_B[5],mul_res1[4205]);
multi_7x28 multi_7x28_mod_4206(clk,rst,matrix_A[4206],matrix_B[6],mul_res1[4206]);
multi_7x28 multi_7x28_mod_4207(clk,rst,matrix_A[4207],matrix_B[7],mul_res1[4207]);
multi_7x28 multi_7x28_mod_4208(clk,rst,matrix_A[4208],matrix_B[8],mul_res1[4208]);
multi_7x28 multi_7x28_mod_4209(clk,rst,matrix_A[4209],matrix_B[9],mul_res1[4209]);
multi_7x28 multi_7x28_mod_4210(clk,rst,matrix_A[4210],matrix_B[10],mul_res1[4210]);
multi_7x28 multi_7x28_mod_4211(clk,rst,matrix_A[4211],matrix_B[11],mul_res1[4211]);
multi_7x28 multi_7x28_mod_4212(clk,rst,matrix_A[4212],matrix_B[12],mul_res1[4212]);
multi_7x28 multi_7x28_mod_4213(clk,rst,matrix_A[4213],matrix_B[13],mul_res1[4213]);
multi_7x28 multi_7x28_mod_4214(clk,rst,matrix_A[4214],matrix_B[14],mul_res1[4214]);
multi_7x28 multi_7x28_mod_4215(clk,rst,matrix_A[4215],matrix_B[15],mul_res1[4215]);
multi_7x28 multi_7x28_mod_4216(clk,rst,matrix_A[4216],matrix_B[16],mul_res1[4216]);
multi_7x28 multi_7x28_mod_4217(clk,rst,matrix_A[4217],matrix_B[17],mul_res1[4217]);
multi_7x28 multi_7x28_mod_4218(clk,rst,matrix_A[4218],matrix_B[18],mul_res1[4218]);
multi_7x28 multi_7x28_mod_4219(clk,rst,matrix_A[4219],matrix_B[19],mul_res1[4219]);
multi_7x28 multi_7x28_mod_4220(clk,rst,matrix_A[4220],matrix_B[20],mul_res1[4220]);
multi_7x28 multi_7x28_mod_4221(clk,rst,matrix_A[4221],matrix_B[21],mul_res1[4221]);
multi_7x28 multi_7x28_mod_4222(clk,rst,matrix_A[4222],matrix_B[22],mul_res1[4222]);
multi_7x28 multi_7x28_mod_4223(clk,rst,matrix_A[4223],matrix_B[23],mul_res1[4223]);
multi_7x28 multi_7x28_mod_4224(clk,rst,matrix_A[4224],matrix_B[24],mul_res1[4224]);
multi_7x28 multi_7x28_mod_4225(clk,rst,matrix_A[4225],matrix_B[25],mul_res1[4225]);
multi_7x28 multi_7x28_mod_4226(clk,rst,matrix_A[4226],matrix_B[26],mul_res1[4226]);
multi_7x28 multi_7x28_mod_4227(clk,rst,matrix_A[4227],matrix_B[27],mul_res1[4227]);
multi_7x28 multi_7x28_mod_4228(clk,rst,matrix_A[4228],matrix_B[28],mul_res1[4228]);
multi_7x28 multi_7x28_mod_4229(clk,rst,matrix_A[4229],matrix_B[29],mul_res1[4229]);
multi_7x28 multi_7x28_mod_4230(clk,rst,matrix_A[4230],matrix_B[30],mul_res1[4230]);
multi_7x28 multi_7x28_mod_4231(clk,rst,matrix_A[4231],matrix_B[31],mul_res1[4231]);
multi_7x28 multi_7x28_mod_4232(clk,rst,matrix_A[4232],matrix_B[32],mul_res1[4232]);
multi_7x28 multi_7x28_mod_4233(clk,rst,matrix_A[4233],matrix_B[33],mul_res1[4233]);
multi_7x28 multi_7x28_mod_4234(clk,rst,matrix_A[4234],matrix_B[34],mul_res1[4234]);
multi_7x28 multi_7x28_mod_4235(clk,rst,matrix_A[4235],matrix_B[35],mul_res1[4235]);
multi_7x28 multi_7x28_mod_4236(clk,rst,matrix_A[4236],matrix_B[36],mul_res1[4236]);
multi_7x28 multi_7x28_mod_4237(clk,rst,matrix_A[4237],matrix_B[37],mul_res1[4237]);
multi_7x28 multi_7x28_mod_4238(clk,rst,matrix_A[4238],matrix_B[38],mul_res1[4238]);
multi_7x28 multi_7x28_mod_4239(clk,rst,matrix_A[4239],matrix_B[39],mul_res1[4239]);
multi_7x28 multi_7x28_mod_4240(clk,rst,matrix_A[4240],matrix_B[40],mul_res1[4240]);
multi_7x28 multi_7x28_mod_4241(clk,rst,matrix_A[4241],matrix_B[41],mul_res1[4241]);
multi_7x28 multi_7x28_mod_4242(clk,rst,matrix_A[4242],matrix_B[42],mul_res1[4242]);
multi_7x28 multi_7x28_mod_4243(clk,rst,matrix_A[4243],matrix_B[43],mul_res1[4243]);
multi_7x28 multi_7x28_mod_4244(clk,rst,matrix_A[4244],matrix_B[44],mul_res1[4244]);
multi_7x28 multi_7x28_mod_4245(clk,rst,matrix_A[4245],matrix_B[45],mul_res1[4245]);
multi_7x28 multi_7x28_mod_4246(clk,rst,matrix_A[4246],matrix_B[46],mul_res1[4246]);
multi_7x28 multi_7x28_mod_4247(clk,rst,matrix_A[4247],matrix_B[47],mul_res1[4247]);
multi_7x28 multi_7x28_mod_4248(clk,rst,matrix_A[4248],matrix_B[48],mul_res1[4248]);
multi_7x28 multi_7x28_mod_4249(clk,rst,matrix_A[4249],matrix_B[49],mul_res1[4249]);
multi_7x28 multi_7x28_mod_4250(clk,rst,matrix_A[4250],matrix_B[50],mul_res1[4250]);
multi_7x28 multi_7x28_mod_4251(clk,rst,matrix_A[4251],matrix_B[51],mul_res1[4251]);
multi_7x28 multi_7x28_mod_4252(clk,rst,matrix_A[4252],matrix_B[52],mul_res1[4252]);
multi_7x28 multi_7x28_mod_4253(clk,rst,matrix_A[4253],matrix_B[53],mul_res1[4253]);
multi_7x28 multi_7x28_mod_4254(clk,rst,matrix_A[4254],matrix_B[54],mul_res1[4254]);
multi_7x28 multi_7x28_mod_4255(clk,rst,matrix_A[4255],matrix_B[55],mul_res1[4255]);
multi_7x28 multi_7x28_mod_4256(clk,rst,matrix_A[4256],matrix_B[56],mul_res1[4256]);
multi_7x28 multi_7x28_mod_4257(clk,rst,matrix_A[4257],matrix_B[57],mul_res1[4257]);
multi_7x28 multi_7x28_mod_4258(clk,rst,matrix_A[4258],matrix_B[58],mul_res1[4258]);
multi_7x28 multi_7x28_mod_4259(clk,rst,matrix_A[4259],matrix_B[59],mul_res1[4259]);
multi_7x28 multi_7x28_mod_4260(clk,rst,matrix_A[4260],matrix_B[60],mul_res1[4260]);
multi_7x28 multi_7x28_mod_4261(clk,rst,matrix_A[4261],matrix_B[61],mul_res1[4261]);
multi_7x28 multi_7x28_mod_4262(clk,rst,matrix_A[4262],matrix_B[62],mul_res1[4262]);
multi_7x28 multi_7x28_mod_4263(clk,rst,matrix_A[4263],matrix_B[63],mul_res1[4263]);
multi_7x28 multi_7x28_mod_4264(clk,rst,matrix_A[4264],matrix_B[64],mul_res1[4264]);
multi_7x28 multi_7x28_mod_4265(clk,rst,matrix_A[4265],matrix_B[65],mul_res1[4265]);
multi_7x28 multi_7x28_mod_4266(clk,rst,matrix_A[4266],matrix_B[66],mul_res1[4266]);
multi_7x28 multi_7x28_mod_4267(clk,rst,matrix_A[4267],matrix_B[67],mul_res1[4267]);
multi_7x28 multi_7x28_mod_4268(clk,rst,matrix_A[4268],matrix_B[68],mul_res1[4268]);
multi_7x28 multi_7x28_mod_4269(clk,rst,matrix_A[4269],matrix_B[69],mul_res1[4269]);
multi_7x28 multi_7x28_mod_4270(clk,rst,matrix_A[4270],matrix_B[70],mul_res1[4270]);
multi_7x28 multi_7x28_mod_4271(clk,rst,matrix_A[4271],matrix_B[71],mul_res1[4271]);
multi_7x28 multi_7x28_mod_4272(clk,rst,matrix_A[4272],matrix_B[72],mul_res1[4272]);
multi_7x28 multi_7x28_mod_4273(clk,rst,matrix_A[4273],matrix_B[73],mul_res1[4273]);
multi_7x28 multi_7x28_mod_4274(clk,rst,matrix_A[4274],matrix_B[74],mul_res1[4274]);
multi_7x28 multi_7x28_mod_4275(clk,rst,matrix_A[4275],matrix_B[75],mul_res1[4275]);
multi_7x28 multi_7x28_mod_4276(clk,rst,matrix_A[4276],matrix_B[76],mul_res1[4276]);
multi_7x28 multi_7x28_mod_4277(clk,rst,matrix_A[4277],matrix_B[77],mul_res1[4277]);
multi_7x28 multi_7x28_mod_4278(clk,rst,matrix_A[4278],matrix_B[78],mul_res1[4278]);
multi_7x28 multi_7x28_mod_4279(clk,rst,matrix_A[4279],matrix_B[79],mul_res1[4279]);
multi_7x28 multi_7x28_mod_4280(clk,rst,matrix_A[4280],matrix_B[80],mul_res1[4280]);
multi_7x28 multi_7x28_mod_4281(clk,rst,matrix_A[4281],matrix_B[81],mul_res1[4281]);
multi_7x28 multi_7x28_mod_4282(clk,rst,matrix_A[4282],matrix_B[82],mul_res1[4282]);
multi_7x28 multi_7x28_mod_4283(clk,rst,matrix_A[4283],matrix_B[83],mul_res1[4283]);
multi_7x28 multi_7x28_mod_4284(clk,rst,matrix_A[4284],matrix_B[84],mul_res1[4284]);
multi_7x28 multi_7x28_mod_4285(clk,rst,matrix_A[4285],matrix_B[85],mul_res1[4285]);
multi_7x28 multi_7x28_mod_4286(clk,rst,matrix_A[4286],matrix_B[86],mul_res1[4286]);
multi_7x28 multi_7x28_mod_4287(clk,rst,matrix_A[4287],matrix_B[87],mul_res1[4287]);
multi_7x28 multi_7x28_mod_4288(clk,rst,matrix_A[4288],matrix_B[88],mul_res1[4288]);
multi_7x28 multi_7x28_mod_4289(clk,rst,matrix_A[4289],matrix_B[89],mul_res1[4289]);
multi_7x28 multi_7x28_mod_4290(clk,rst,matrix_A[4290],matrix_B[90],mul_res1[4290]);
multi_7x28 multi_7x28_mod_4291(clk,rst,matrix_A[4291],matrix_B[91],mul_res1[4291]);
multi_7x28 multi_7x28_mod_4292(clk,rst,matrix_A[4292],matrix_B[92],mul_res1[4292]);
multi_7x28 multi_7x28_mod_4293(clk,rst,matrix_A[4293],matrix_B[93],mul_res1[4293]);
multi_7x28 multi_7x28_mod_4294(clk,rst,matrix_A[4294],matrix_B[94],mul_res1[4294]);
multi_7x28 multi_7x28_mod_4295(clk,rst,matrix_A[4295],matrix_B[95],mul_res1[4295]);
multi_7x28 multi_7x28_mod_4296(clk,rst,matrix_A[4296],matrix_B[96],mul_res1[4296]);
multi_7x28 multi_7x28_mod_4297(clk,rst,matrix_A[4297],matrix_B[97],mul_res1[4297]);
multi_7x28 multi_7x28_mod_4298(clk,rst,matrix_A[4298],matrix_B[98],mul_res1[4298]);
multi_7x28 multi_7x28_mod_4299(clk,rst,matrix_A[4299],matrix_B[99],mul_res1[4299]);
multi_7x28 multi_7x28_mod_4300(clk,rst,matrix_A[4300],matrix_B[100],mul_res1[4300]);
multi_7x28 multi_7x28_mod_4301(clk,rst,matrix_A[4301],matrix_B[101],mul_res1[4301]);
multi_7x28 multi_7x28_mod_4302(clk,rst,matrix_A[4302],matrix_B[102],mul_res1[4302]);
multi_7x28 multi_7x28_mod_4303(clk,rst,matrix_A[4303],matrix_B[103],mul_res1[4303]);
multi_7x28 multi_7x28_mod_4304(clk,rst,matrix_A[4304],matrix_B[104],mul_res1[4304]);
multi_7x28 multi_7x28_mod_4305(clk,rst,matrix_A[4305],matrix_B[105],mul_res1[4305]);
multi_7x28 multi_7x28_mod_4306(clk,rst,matrix_A[4306],matrix_B[106],mul_res1[4306]);
multi_7x28 multi_7x28_mod_4307(clk,rst,matrix_A[4307],matrix_B[107],mul_res1[4307]);
multi_7x28 multi_7x28_mod_4308(clk,rst,matrix_A[4308],matrix_B[108],mul_res1[4308]);
multi_7x28 multi_7x28_mod_4309(clk,rst,matrix_A[4309],matrix_B[109],mul_res1[4309]);
multi_7x28 multi_7x28_mod_4310(clk,rst,matrix_A[4310],matrix_B[110],mul_res1[4310]);
multi_7x28 multi_7x28_mod_4311(clk,rst,matrix_A[4311],matrix_B[111],mul_res1[4311]);
multi_7x28 multi_7x28_mod_4312(clk,rst,matrix_A[4312],matrix_B[112],mul_res1[4312]);
multi_7x28 multi_7x28_mod_4313(clk,rst,matrix_A[4313],matrix_B[113],mul_res1[4313]);
multi_7x28 multi_7x28_mod_4314(clk,rst,matrix_A[4314],matrix_B[114],mul_res1[4314]);
multi_7x28 multi_7x28_mod_4315(clk,rst,matrix_A[4315],matrix_B[115],mul_res1[4315]);
multi_7x28 multi_7x28_mod_4316(clk,rst,matrix_A[4316],matrix_B[116],mul_res1[4316]);
multi_7x28 multi_7x28_mod_4317(clk,rst,matrix_A[4317],matrix_B[117],mul_res1[4317]);
multi_7x28 multi_7x28_mod_4318(clk,rst,matrix_A[4318],matrix_B[118],mul_res1[4318]);
multi_7x28 multi_7x28_mod_4319(clk,rst,matrix_A[4319],matrix_B[119],mul_res1[4319]);
multi_7x28 multi_7x28_mod_4320(clk,rst,matrix_A[4320],matrix_B[120],mul_res1[4320]);
multi_7x28 multi_7x28_mod_4321(clk,rst,matrix_A[4321],matrix_B[121],mul_res1[4321]);
multi_7x28 multi_7x28_mod_4322(clk,rst,matrix_A[4322],matrix_B[122],mul_res1[4322]);
multi_7x28 multi_7x28_mod_4323(clk,rst,matrix_A[4323],matrix_B[123],mul_res1[4323]);
multi_7x28 multi_7x28_mod_4324(clk,rst,matrix_A[4324],matrix_B[124],mul_res1[4324]);
multi_7x28 multi_7x28_mod_4325(clk,rst,matrix_A[4325],matrix_B[125],mul_res1[4325]);
multi_7x28 multi_7x28_mod_4326(clk,rst,matrix_A[4326],matrix_B[126],mul_res1[4326]);
multi_7x28 multi_7x28_mod_4327(clk,rst,matrix_A[4327],matrix_B[127],mul_res1[4327]);
multi_7x28 multi_7x28_mod_4328(clk,rst,matrix_A[4328],matrix_B[128],mul_res1[4328]);
multi_7x28 multi_7x28_mod_4329(clk,rst,matrix_A[4329],matrix_B[129],mul_res1[4329]);
multi_7x28 multi_7x28_mod_4330(clk,rst,matrix_A[4330],matrix_B[130],mul_res1[4330]);
multi_7x28 multi_7x28_mod_4331(clk,rst,matrix_A[4331],matrix_B[131],mul_res1[4331]);
multi_7x28 multi_7x28_mod_4332(clk,rst,matrix_A[4332],matrix_B[132],mul_res1[4332]);
multi_7x28 multi_7x28_mod_4333(clk,rst,matrix_A[4333],matrix_B[133],mul_res1[4333]);
multi_7x28 multi_7x28_mod_4334(clk,rst,matrix_A[4334],matrix_B[134],mul_res1[4334]);
multi_7x28 multi_7x28_mod_4335(clk,rst,matrix_A[4335],matrix_B[135],mul_res1[4335]);
multi_7x28 multi_7x28_mod_4336(clk,rst,matrix_A[4336],matrix_B[136],mul_res1[4336]);
multi_7x28 multi_7x28_mod_4337(clk,rst,matrix_A[4337],matrix_B[137],mul_res1[4337]);
multi_7x28 multi_7x28_mod_4338(clk,rst,matrix_A[4338],matrix_B[138],mul_res1[4338]);
multi_7x28 multi_7x28_mod_4339(clk,rst,matrix_A[4339],matrix_B[139],mul_res1[4339]);
multi_7x28 multi_7x28_mod_4340(clk,rst,matrix_A[4340],matrix_B[140],mul_res1[4340]);
multi_7x28 multi_7x28_mod_4341(clk,rst,matrix_A[4341],matrix_B[141],mul_res1[4341]);
multi_7x28 multi_7x28_mod_4342(clk,rst,matrix_A[4342],matrix_B[142],mul_res1[4342]);
multi_7x28 multi_7x28_mod_4343(clk,rst,matrix_A[4343],matrix_B[143],mul_res1[4343]);
multi_7x28 multi_7x28_mod_4344(clk,rst,matrix_A[4344],matrix_B[144],mul_res1[4344]);
multi_7x28 multi_7x28_mod_4345(clk,rst,matrix_A[4345],matrix_B[145],mul_res1[4345]);
multi_7x28 multi_7x28_mod_4346(clk,rst,matrix_A[4346],matrix_B[146],mul_res1[4346]);
multi_7x28 multi_7x28_mod_4347(clk,rst,matrix_A[4347],matrix_B[147],mul_res1[4347]);
multi_7x28 multi_7x28_mod_4348(clk,rst,matrix_A[4348],matrix_B[148],mul_res1[4348]);
multi_7x28 multi_7x28_mod_4349(clk,rst,matrix_A[4349],matrix_B[149],mul_res1[4349]);
multi_7x28 multi_7x28_mod_4350(clk,rst,matrix_A[4350],matrix_B[150],mul_res1[4350]);
multi_7x28 multi_7x28_mod_4351(clk,rst,matrix_A[4351],matrix_B[151],mul_res1[4351]);
multi_7x28 multi_7x28_mod_4352(clk,rst,matrix_A[4352],matrix_B[152],mul_res1[4352]);
multi_7x28 multi_7x28_mod_4353(clk,rst,matrix_A[4353],matrix_B[153],mul_res1[4353]);
multi_7x28 multi_7x28_mod_4354(clk,rst,matrix_A[4354],matrix_B[154],mul_res1[4354]);
multi_7x28 multi_7x28_mod_4355(clk,rst,matrix_A[4355],matrix_B[155],mul_res1[4355]);
multi_7x28 multi_7x28_mod_4356(clk,rst,matrix_A[4356],matrix_B[156],mul_res1[4356]);
multi_7x28 multi_7x28_mod_4357(clk,rst,matrix_A[4357],matrix_B[157],mul_res1[4357]);
multi_7x28 multi_7x28_mod_4358(clk,rst,matrix_A[4358],matrix_B[158],mul_res1[4358]);
multi_7x28 multi_7x28_mod_4359(clk,rst,matrix_A[4359],matrix_B[159],mul_res1[4359]);
multi_7x28 multi_7x28_mod_4360(clk,rst,matrix_A[4360],matrix_B[160],mul_res1[4360]);
multi_7x28 multi_7x28_mod_4361(clk,rst,matrix_A[4361],matrix_B[161],mul_res1[4361]);
multi_7x28 multi_7x28_mod_4362(clk,rst,matrix_A[4362],matrix_B[162],mul_res1[4362]);
multi_7x28 multi_7x28_mod_4363(clk,rst,matrix_A[4363],matrix_B[163],mul_res1[4363]);
multi_7x28 multi_7x28_mod_4364(clk,rst,matrix_A[4364],matrix_B[164],mul_res1[4364]);
multi_7x28 multi_7x28_mod_4365(clk,rst,matrix_A[4365],matrix_B[165],mul_res1[4365]);
multi_7x28 multi_7x28_mod_4366(clk,rst,matrix_A[4366],matrix_B[166],mul_res1[4366]);
multi_7x28 multi_7x28_mod_4367(clk,rst,matrix_A[4367],matrix_B[167],mul_res1[4367]);
multi_7x28 multi_7x28_mod_4368(clk,rst,matrix_A[4368],matrix_B[168],mul_res1[4368]);
multi_7x28 multi_7x28_mod_4369(clk,rst,matrix_A[4369],matrix_B[169],mul_res1[4369]);
multi_7x28 multi_7x28_mod_4370(clk,rst,matrix_A[4370],matrix_B[170],mul_res1[4370]);
multi_7x28 multi_7x28_mod_4371(clk,rst,matrix_A[4371],matrix_B[171],mul_res1[4371]);
multi_7x28 multi_7x28_mod_4372(clk,rst,matrix_A[4372],matrix_B[172],mul_res1[4372]);
multi_7x28 multi_7x28_mod_4373(clk,rst,matrix_A[4373],matrix_B[173],mul_res1[4373]);
multi_7x28 multi_7x28_mod_4374(clk,rst,matrix_A[4374],matrix_B[174],mul_res1[4374]);
multi_7x28 multi_7x28_mod_4375(clk,rst,matrix_A[4375],matrix_B[175],mul_res1[4375]);
multi_7x28 multi_7x28_mod_4376(clk,rst,matrix_A[4376],matrix_B[176],mul_res1[4376]);
multi_7x28 multi_7x28_mod_4377(clk,rst,matrix_A[4377],matrix_B[177],mul_res1[4377]);
multi_7x28 multi_7x28_mod_4378(clk,rst,matrix_A[4378],matrix_B[178],mul_res1[4378]);
multi_7x28 multi_7x28_mod_4379(clk,rst,matrix_A[4379],matrix_B[179],mul_res1[4379]);
multi_7x28 multi_7x28_mod_4380(clk,rst,matrix_A[4380],matrix_B[180],mul_res1[4380]);
multi_7x28 multi_7x28_mod_4381(clk,rst,matrix_A[4381],matrix_B[181],mul_res1[4381]);
multi_7x28 multi_7x28_mod_4382(clk,rst,matrix_A[4382],matrix_B[182],mul_res1[4382]);
multi_7x28 multi_7x28_mod_4383(clk,rst,matrix_A[4383],matrix_B[183],mul_res1[4383]);
multi_7x28 multi_7x28_mod_4384(clk,rst,matrix_A[4384],matrix_B[184],mul_res1[4384]);
multi_7x28 multi_7x28_mod_4385(clk,rst,matrix_A[4385],matrix_B[185],mul_res1[4385]);
multi_7x28 multi_7x28_mod_4386(clk,rst,matrix_A[4386],matrix_B[186],mul_res1[4386]);
multi_7x28 multi_7x28_mod_4387(clk,rst,matrix_A[4387],matrix_B[187],mul_res1[4387]);
multi_7x28 multi_7x28_mod_4388(clk,rst,matrix_A[4388],matrix_B[188],mul_res1[4388]);
multi_7x28 multi_7x28_mod_4389(clk,rst,matrix_A[4389],matrix_B[189],mul_res1[4389]);
multi_7x28 multi_7x28_mod_4390(clk,rst,matrix_A[4390],matrix_B[190],mul_res1[4390]);
multi_7x28 multi_7x28_mod_4391(clk,rst,matrix_A[4391],matrix_B[191],mul_res1[4391]);
multi_7x28 multi_7x28_mod_4392(clk,rst,matrix_A[4392],matrix_B[192],mul_res1[4392]);
multi_7x28 multi_7x28_mod_4393(clk,rst,matrix_A[4393],matrix_B[193],mul_res1[4393]);
multi_7x28 multi_7x28_mod_4394(clk,rst,matrix_A[4394],matrix_B[194],mul_res1[4394]);
multi_7x28 multi_7x28_mod_4395(clk,rst,matrix_A[4395],matrix_B[195],mul_res1[4395]);
multi_7x28 multi_7x28_mod_4396(clk,rst,matrix_A[4396],matrix_B[196],mul_res1[4396]);
multi_7x28 multi_7x28_mod_4397(clk,rst,matrix_A[4397],matrix_B[197],mul_res1[4397]);
multi_7x28 multi_7x28_mod_4398(clk,rst,matrix_A[4398],matrix_B[198],mul_res1[4398]);
multi_7x28 multi_7x28_mod_4399(clk,rst,matrix_A[4399],matrix_B[199],mul_res1[4399]);
multi_7x28 multi_7x28_mod_4400(clk,rst,matrix_A[4400],matrix_B[0],mul_res1[4400]);
multi_7x28 multi_7x28_mod_4401(clk,rst,matrix_A[4401],matrix_B[1],mul_res1[4401]);
multi_7x28 multi_7x28_mod_4402(clk,rst,matrix_A[4402],matrix_B[2],mul_res1[4402]);
multi_7x28 multi_7x28_mod_4403(clk,rst,matrix_A[4403],matrix_B[3],mul_res1[4403]);
multi_7x28 multi_7x28_mod_4404(clk,rst,matrix_A[4404],matrix_B[4],mul_res1[4404]);
multi_7x28 multi_7x28_mod_4405(clk,rst,matrix_A[4405],matrix_B[5],mul_res1[4405]);
multi_7x28 multi_7x28_mod_4406(clk,rst,matrix_A[4406],matrix_B[6],mul_res1[4406]);
multi_7x28 multi_7x28_mod_4407(clk,rst,matrix_A[4407],matrix_B[7],mul_res1[4407]);
multi_7x28 multi_7x28_mod_4408(clk,rst,matrix_A[4408],matrix_B[8],mul_res1[4408]);
multi_7x28 multi_7x28_mod_4409(clk,rst,matrix_A[4409],matrix_B[9],mul_res1[4409]);
multi_7x28 multi_7x28_mod_4410(clk,rst,matrix_A[4410],matrix_B[10],mul_res1[4410]);
multi_7x28 multi_7x28_mod_4411(clk,rst,matrix_A[4411],matrix_B[11],mul_res1[4411]);
multi_7x28 multi_7x28_mod_4412(clk,rst,matrix_A[4412],matrix_B[12],mul_res1[4412]);
multi_7x28 multi_7x28_mod_4413(clk,rst,matrix_A[4413],matrix_B[13],mul_res1[4413]);
multi_7x28 multi_7x28_mod_4414(clk,rst,matrix_A[4414],matrix_B[14],mul_res1[4414]);
multi_7x28 multi_7x28_mod_4415(clk,rst,matrix_A[4415],matrix_B[15],mul_res1[4415]);
multi_7x28 multi_7x28_mod_4416(clk,rst,matrix_A[4416],matrix_B[16],mul_res1[4416]);
multi_7x28 multi_7x28_mod_4417(clk,rst,matrix_A[4417],matrix_B[17],mul_res1[4417]);
multi_7x28 multi_7x28_mod_4418(clk,rst,matrix_A[4418],matrix_B[18],mul_res1[4418]);
multi_7x28 multi_7x28_mod_4419(clk,rst,matrix_A[4419],matrix_B[19],mul_res1[4419]);
multi_7x28 multi_7x28_mod_4420(clk,rst,matrix_A[4420],matrix_B[20],mul_res1[4420]);
multi_7x28 multi_7x28_mod_4421(clk,rst,matrix_A[4421],matrix_B[21],mul_res1[4421]);
multi_7x28 multi_7x28_mod_4422(clk,rst,matrix_A[4422],matrix_B[22],mul_res1[4422]);
multi_7x28 multi_7x28_mod_4423(clk,rst,matrix_A[4423],matrix_B[23],mul_res1[4423]);
multi_7x28 multi_7x28_mod_4424(clk,rst,matrix_A[4424],matrix_B[24],mul_res1[4424]);
multi_7x28 multi_7x28_mod_4425(clk,rst,matrix_A[4425],matrix_B[25],mul_res1[4425]);
multi_7x28 multi_7x28_mod_4426(clk,rst,matrix_A[4426],matrix_B[26],mul_res1[4426]);
multi_7x28 multi_7x28_mod_4427(clk,rst,matrix_A[4427],matrix_B[27],mul_res1[4427]);
multi_7x28 multi_7x28_mod_4428(clk,rst,matrix_A[4428],matrix_B[28],mul_res1[4428]);
multi_7x28 multi_7x28_mod_4429(clk,rst,matrix_A[4429],matrix_B[29],mul_res1[4429]);
multi_7x28 multi_7x28_mod_4430(clk,rst,matrix_A[4430],matrix_B[30],mul_res1[4430]);
multi_7x28 multi_7x28_mod_4431(clk,rst,matrix_A[4431],matrix_B[31],mul_res1[4431]);
multi_7x28 multi_7x28_mod_4432(clk,rst,matrix_A[4432],matrix_B[32],mul_res1[4432]);
multi_7x28 multi_7x28_mod_4433(clk,rst,matrix_A[4433],matrix_B[33],mul_res1[4433]);
multi_7x28 multi_7x28_mod_4434(clk,rst,matrix_A[4434],matrix_B[34],mul_res1[4434]);
multi_7x28 multi_7x28_mod_4435(clk,rst,matrix_A[4435],matrix_B[35],mul_res1[4435]);
multi_7x28 multi_7x28_mod_4436(clk,rst,matrix_A[4436],matrix_B[36],mul_res1[4436]);
multi_7x28 multi_7x28_mod_4437(clk,rst,matrix_A[4437],matrix_B[37],mul_res1[4437]);
multi_7x28 multi_7x28_mod_4438(clk,rst,matrix_A[4438],matrix_B[38],mul_res1[4438]);
multi_7x28 multi_7x28_mod_4439(clk,rst,matrix_A[4439],matrix_B[39],mul_res1[4439]);
multi_7x28 multi_7x28_mod_4440(clk,rst,matrix_A[4440],matrix_B[40],mul_res1[4440]);
multi_7x28 multi_7x28_mod_4441(clk,rst,matrix_A[4441],matrix_B[41],mul_res1[4441]);
multi_7x28 multi_7x28_mod_4442(clk,rst,matrix_A[4442],matrix_B[42],mul_res1[4442]);
multi_7x28 multi_7x28_mod_4443(clk,rst,matrix_A[4443],matrix_B[43],mul_res1[4443]);
multi_7x28 multi_7x28_mod_4444(clk,rst,matrix_A[4444],matrix_B[44],mul_res1[4444]);
multi_7x28 multi_7x28_mod_4445(clk,rst,matrix_A[4445],matrix_B[45],mul_res1[4445]);
multi_7x28 multi_7x28_mod_4446(clk,rst,matrix_A[4446],matrix_B[46],mul_res1[4446]);
multi_7x28 multi_7x28_mod_4447(clk,rst,matrix_A[4447],matrix_B[47],mul_res1[4447]);
multi_7x28 multi_7x28_mod_4448(clk,rst,matrix_A[4448],matrix_B[48],mul_res1[4448]);
multi_7x28 multi_7x28_mod_4449(clk,rst,matrix_A[4449],matrix_B[49],mul_res1[4449]);
multi_7x28 multi_7x28_mod_4450(clk,rst,matrix_A[4450],matrix_B[50],mul_res1[4450]);
multi_7x28 multi_7x28_mod_4451(clk,rst,matrix_A[4451],matrix_B[51],mul_res1[4451]);
multi_7x28 multi_7x28_mod_4452(clk,rst,matrix_A[4452],matrix_B[52],mul_res1[4452]);
multi_7x28 multi_7x28_mod_4453(clk,rst,matrix_A[4453],matrix_B[53],mul_res1[4453]);
multi_7x28 multi_7x28_mod_4454(clk,rst,matrix_A[4454],matrix_B[54],mul_res1[4454]);
multi_7x28 multi_7x28_mod_4455(clk,rst,matrix_A[4455],matrix_B[55],mul_res1[4455]);
multi_7x28 multi_7x28_mod_4456(clk,rst,matrix_A[4456],matrix_B[56],mul_res1[4456]);
multi_7x28 multi_7x28_mod_4457(clk,rst,matrix_A[4457],matrix_B[57],mul_res1[4457]);
multi_7x28 multi_7x28_mod_4458(clk,rst,matrix_A[4458],matrix_B[58],mul_res1[4458]);
multi_7x28 multi_7x28_mod_4459(clk,rst,matrix_A[4459],matrix_B[59],mul_res1[4459]);
multi_7x28 multi_7x28_mod_4460(clk,rst,matrix_A[4460],matrix_B[60],mul_res1[4460]);
multi_7x28 multi_7x28_mod_4461(clk,rst,matrix_A[4461],matrix_B[61],mul_res1[4461]);
multi_7x28 multi_7x28_mod_4462(clk,rst,matrix_A[4462],matrix_B[62],mul_res1[4462]);
multi_7x28 multi_7x28_mod_4463(clk,rst,matrix_A[4463],matrix_B[63],mul_res1[4463]);
multi_7x28 multi_7x28_mod_4464(clk,rst,matrix_A[4464],matrix_B[64],mul_res1[4464]);
multi_7x28 multi_7x28_mod_4465(clk,rst,matrix_A[4465],matrix_B[65],mul_res1[4465]);
multi_7x28 multi_7x28_mod_4466(clk,rst,matrix_A[4466],matrix_B[66],mul_res1[4466]);
multi_7x28 multi_7x28_mod_4467(clk,rst,matrix_A[4467],matrix_B[67],mul_res1[4467]);
multi_7x28 multi_7x28_mod_4468(clk,rst,matrix_A[4468],matrix_B[68],mul_res1[4468]);
multi_7x28 multi_7x28_mod_4469(clk,rst,matrix_A[4469],matrix_B[69],mul_res1[4469]);
multi_7x28 multi_7x28_mod_4470(clk,rst,matrix_A[4470],matrix_B[70],mul_res1[4470]);
multi_7x28 multi_7x28_mod_4471(clk,rst,matrix_A[4471],matrix_B[71],mul_res1[4471]);
multi_7x28 multi_7x28_mod_4472(clk,rst,matrix_A[4472],matrix_B[72],mul_res1[4472]);
multi_7x28 multi_7x28_mod_4473(clk,rst,matrix_A[4473],matrix_B[73],mul_res1[4473]);
multi_7x28 multi_7x28_mod_4474(clk,rst,matrix_A[4474],matrix_B[74],mul_res1[4474]);
multi_7x28 multi_7x28_mod_4475(clk,rst,matrix_A[4475],matrix_B[75],mul_res1[4475]);
multi_7x28 multi_7x28_mod_4476(clk,rst,matrix_A[4476],matrix_B[76],mul_res1[4476]);
multi_7x28 multi_7x28_mod_4477(clk,rst,matrix_A[4477],matrix_B[77],mul_res1[4477]);
multi_7x28 multi_7x28_mod_4478(clk,rst,matrix_A[4478],matrix_B[78],mul_res1[4478]);
multi_7x28 multi_7x28_mod_4479(clk,rst,matrix_A[4479],matrix_B[79],mul_res1[4479]);
multi_7x28 multi_7x28_mod_4480(clk,rst,matrix_A[4480],matrix_B[80],mul_res1[4480]);
multi_7x28 multi_7x28_mod_4481(clk,rst,matrix_A[4481],matrix_B[81],mul_res1[4481]);
multi_7x28 multi_7x28_mod_4482(clk,rst,matrix_A[4482],matrix_B[82],mul_res1[4482]);
multi_7x28 multi_7x28_mod_4483(clk,rst,matrix_A[4483],matrix_B[83],mul_res1[4483]);
multi_7x28 multi_7x28_mod_4484(clk,rst,matrix_A[4484],matrix_B[84],mul_res1[4484]);
multi_7x28 multi_7x28_mod_4485(clk,rst,matrix_A[4485],matrix_B[85],mul_res1[4485]);
multi_7x28 multi_7x28_mod_4486(clk,rst,matrix_A[4486],matrix_B[86],mul_res1[4486]);
multi_7x28 multi_7x28_mod_4487(clk,rst,matrix_A[4487],matrix_B[87],mul_res1[4487]);
multi_7x28 multi_7x28_mod_4488(clk,rst,matrix_A[4488],matrix_B[88],mul_res1[4488]);
multi_7x28 multi_7x28_mod_4489(clk,rst,matrix_A[4489],matrix_B[89],mul_res1[4489]);
multi_7x28 multi_7x28_mod_4490(clk,rst,matrix_A[4490],matrix_B[90],mul_res1[4490]);
multi_7x28 multi_7x28_mod_4491(clk,rst,matrix_A[4491],matrix_B[91],mul_res1[4491]);
multi_7x28 multi_7x28_mod_4492(clk,rst,matrix_A[4492],matrix_B[92],mul_res1[4492]);
multi_7x28 multi_7x28_mod_4493(clk,rst,matrix_A[4493],matrix_B[93],mul_res1[4493]);
multi_7x28 multi_7x28_mod_4494(clk,rst,matrix_A[4494],matrix_B[94],mul_res1[4494]);
multi_7x28 multi_7x28_mod_4495(clk,rst,matrix_A[4495],matrix_B[95],mul_res1[4495]);
multi_7x28 multi_7x28_mod_4496(clk,rst,matrix_A[4496],matrix_B[96],mul_res1[4496]);
multi_7x28 multi_7x28_mod_4497(clk,rst,matrix_A[4497],matrix_B[97],mul_res1[4497]);
multi_7x28 multi_7x28_mod_4498(clk,rst,matrix_A[4498],matrix_B[98],mul_res1[4498]);
multi_7x28 multi_7x28_mod_4499(clk,rst,matrix_A[4499],matrix_B[99],mul_res1[4499]);
multi_7x28 multi_7x28_mod_4500(clk,rst,matrix_A[4500],matrix_B[100],mul_res1[4500]);
multi_7x28 multi_7x28_mod_4501(clk,rst,matrix_A[4501],matrix_B[101],mul_res1[4501]);
multi_7x28 multi_7x28_mod_4502(clk,rst,matrix_A[4502],matrix_B[102],mul_res1[4502]);
multi_7x28 multi_7x28_mod_4503(clk,rst,matrix_A[4503],matrix_B[103],mul_res1[4503]);
multi_7x28 multi_7x28_mod_4504(clk,rst,matrix_A[4504],matrix_B[104],mul_res1[4504]);
multi_7x28 multi_7x28_mod_4505(clk,rst,matrix_A[4505],matrix_B[105],mul_res1[4505]);
multi_7x28 multi_7x28_mod_4506(clk,rst,matrix_A[4506],matrix_B[106],mul_res1[4506]);
multi_7x28 multi_7x28_mod_4507(clk,rst,matrix_A[4507],matrix_B[107],mul_res1[4507]);
multi_7x28 multi_7x28_mod_4508(clk,rst,matrix_A[4508],matrix_B[108],mul_res1[4508]);
multi_7x28 multi_7x28_mod_4509(clk,rst,matrix_A[4509],matrix_B[109],mul_res1[4509]);
multi_7x28 multi_7x28_mod_4510(clk,rst,matrix_A[4510],matrix_B[110],mul_res1[4510]);
multi_7x28 multi_7x28_mod_4511(clk,rst,matrix_A[4511],matrix_B[111],mul_res1[4511]);
multi_7x28 multi_7x28_mod_4512(clk,rst,matrix_A[4512],matrix_B[112],mul_res1[4512]);
multi_7x28 multi_7x28_mod_4513(clk,rst,matrix_A[4513],matrix_B[113],mul_res1[4513]);
multi_7x28 multi_7x28_mod_4514(clk,rst,matrix_A[4514],matrix_B[114],mul_res1[4514]);
multi_7x28 multi_7x28_mod_4515(clk,rst,matrix_A[4515],matrix_B[115],mul_res1[4515]);
multi_7x28 multi_7x28_mod_4516(clk,rst,matrix_A[4516],matrix_B[116],mul_res1[4516]);
multi_7x28 multi_7x28_mod_4517(clk,rst,matrix_A[4517],matrix_B[117],mul_res1[4517]);
multi_7x28 multi_7x28_mod_4518(clk,rst,matrix_A[4518],matrix_B[118],mul_res1[4518]);
multi_7x28 multi_7x28_mod_4519(clk,rst,matrix_A[4519],matrix_B[119],mul_res1[4519]);
multi_7x28 multi_7x28_mod_4520(clk,rst,matrix_A[4520],matrix_B[120],mul_res1[4520]);
multi_7x28 multi_7x28_mod_4521(clk,rst,matrix_A[4521],matrix_B[121],mul_res1[4521]);
multi_7x28 multi_7x28_mod_4522(clk,rst,matrix_A[4522],matrix_B[122],mul_res1[4522]);
multi_7x28 multi_7x28_mod_4523(clk,rst,matrix_A[4523],matrix_B[123],mul_res1[4523]);
multi_7x28 multi_7x28_mod_4524(clk,rst,matrix_A[4524],matrix_B[124],mul_res1[4524]);
multi_7x28 multi_7x28_mod_4525(clk,rst,matrix_A[4525],matrix_B[125],mul_res1[4525]);
multi_7x28 multi_7x28_mod_4526(clk,rst,matrix_A[4526],matrix_B[126],mul_res1[4526]);
multi_7x28 multi_7x28_mod_4527(clk,rst,matrix_A[4527],matrix_B[127],mul_res1[4527]);
multi_7x28 multi_7x28_mod_4528(clk,rst,matrix_A[4528],matrix_B[128],mul_res1[4528]);
multi_7x28 multi_7x28_mod_4529(clk,rst,matrix_A[4529],matrix_B[129],mul_res1[4529]);
multi_7x28 multi_7x28_mod_4530(clk,rst,matrix_A[4530],matrix_B[130],mul_res1[4530]);
multi_7x28 multi_7x28_mod_4531(clk,rst,matrix_A[4531],matrix_B[131],mul_res1[4531]);
multi_7x28 multi_7x28_mod_4532(clk,rst,matrix_A[4532],matrix_B[132],mul_res1[4532]);
multi_7x28 multi_7x28_mod_4533(clk,rst,matrix_A[4533],matrix_B[133],mul_res1[4533]);
multi_7x28 multi_7x28_mod_4534(clk,rst,matrix_A[4534],matrix_B[134],mul_res1[4534]);
multi_7x28 multi_7x28_mod_4535(clk,rst,matrix_A[4535],matrix_B[135],mul_res1[4535]);
multi_7x28 multi_7x28_mod_4536(clk,rst,matrix_A[4536],matrix_B[136],mul_res1[4536]);
multi_7x28 multi_7x28_mod_4537(clk,rst,matrix_A[4537],matrix_B[137],mul_res1[4537]);
multi_7x28 multi_7x28_mod_4538(clk,rst,matrix_A[4538],matrix_B[138],mul_res1[4538]);
multi_7x28 multi_7x28_mod_4539(clk,rst,matrix_A[4539],matrix_B[139],mul_res1[4539]);
multi_7x28 multi_7x28_mod_4540(clk,rst,matrix_A[4540],matrix_B[140],mul_res1[4540]);
multi_7x28 multi_7x28_mod_4541(clk,rst,matrix_A[4541],matrix_B[141],mul_res1[4541]);
multi_7x28 multi_7x28_mod_4542(clk,rst,matrix_A[4542],matrix_B[142],mul_res1[4542]);
multi_7x28 multi_7x28_mod_4543(clk,rst,matrix_A[4543],matrix_B[143],mul_res1[4543]);
multi_7x28 multi_7x28_mod_4544(clk,rst,matrix_A[4544],matrix_B[144],mul_res1[4544]);
multi_7x28 multi_7x28_mod_4545(clk,rst,matrix_A[4545],matrix_B[145],mul_res1[4545]);
multi_7x28 multi_7x28_mod_4546(clk,rst,matrix_A[4546],matrix_B[146],mul_res1[4546]);
multi_7x28 multi_7x28_mod_4547(clk,rst,matrix_A[4547],matrix_B[147],mul_res1[4547]);
multi_7x28 multi_7x28_mod_4548(clk,rst,matrix_A[4548],matrix_B[148],mul_res1[4548]);
multi_7x28 multi_7x28_mod_4549(clk,rst,matrix_A[4549],matrix_B[149],mul_res1[4549]);
multi_7x28 multi_7x28_mod_4550(clk,rst,matrix_A[4550],matrix_B[150],mul_res1[4550]);
multi_7x28 multi_7x28_mod_4551(clk,rst,matrix_A[4551],matrix_B[151],mul_res1[4551]);
multi_7x28 multi_7x28_mod_4552(clk,rst,matrix_A[4552],matrix_B[152],mul_res1[4552]);
multi_7x28 multi_7x28_mod_4553(clk,rst,matrix_A[4553],matrix_B[153],mul_res1[4553]);
multi_7x28 multi_7x28_mod_4554(clk,rst,matrix_A[4554],matrix_B[154],mul_res1[4554]);
multi_7x28 multi_7x28_mod_4555(clk,rst,matrix_A[4555],matrix_B[155],mul_res1[4555]);
multi_7x28 multi_7x28_mod_4556(clk,rst,matrix_A[4556],matrix_B[156],mul_res1[4556]);
multi_7x28 multi_7x28_mod_4557(clk,rst,matrix_A[4557],matrix_B[157],mul_res1[4557]);
multi_7x28 multi_7x28_mod_4558(clk,rst,matrix_A[4558],matrix_B[158],mul_res1[4558]);
multi_7x28 multi_7x28_mod_4559(clk,rst,matrix_A[4559],matrix_B[159],mul_res1[4559]);
multi_7x28 multi_7x28_mod_4560(clk,rst,matrix_A[4560],matrix_B[160],mul_res1[4560]);
multi_7x28 multi_7x28_mod_4561(clk,rst,matrix_A[4561],matrix_B[161],mul_res1[4561]);
multi_7x28 multi_7x28_mod_4562(clk,rst,matrix_A[4562],matrix_B[162],mul_res1[4562]);
multi_7x28 multi_7x28_mod_4563(clk,rst,matrix_A[4563],matrix_B[163],mul_res1[4563]);
multi_7x28 multi_7x28_mod_4564(clk,rst,matrix_A[4564],matrix_B[164],mul_res1[4564]);
multi_7x28 multi_7x28_mod_4565(clk,rst,matrix_A[4565],matrix_B[165],mul_res1[4565]);
multi_7x28 multi_7x28_mod_4566(clk,rst,matrix_A[4566],matrix_B[166],mul_res1[4566]);
multi_7x28 multi_7x28_mod_4567(clk,rst,matrix_A[4567],matrix_B[167],mul_res1[4567]);
multi_7x28 multi_7x28_mod_4568(clk,rst,matrix_A[4568],matrix_B[168],mul_res1[4568]);
multi_7x28 multi_7x28_mod_4569(clk,rst,matrix_A[4569],matrix_B[169],mul_res1[4569]);
multi_7x28 multi_7x28_mod_4570(clk,rst,matrix_A[4570],matrix_B[170],mul_res1[4570]);
multi_7x28 multi_7x28_mod_4571(clk,rst,matrix_A[4571],matrix_B[171],mul_res1[4571]);
multi_7x28 multi_7x28_mod_4572(clk,rst,matrix_A[4572],matrix_B[172],mul_res1[4572]);
multi_7x28 multi_7x28_mod_4573(clk,rst,matrix_A[4573],matrix_B[173],mul_res1[4573]);
multi_7x28 multi_7x28_mod_4574(clk,rst,matrix_A[4574],matrix_B[174],mul_res1[4574]);
multi_7x28 multi_7x28_mod_4575(clk,rst,matrix_A[4575],matrix_B[175],mul_res1[4575]);
multi_7x28 multi_7x28_mod_4576(clk,rst,matrix_A[4576],matrix_B[176],mul_res1[4576]);
multi_7x28 multi_7x28_mod_4577(clk,rst,matrix_A[4577],matrix_B[177],mul_res1[4577]);
multi_7x28 multi_7x28_mod_4578(clk,rst,matrix_A[4578],matrix_B[178],mul_res1[4578]);
multi_7x28 multi_7x28_mod_4579(clk,rst,matrix_A[4579],matrix_B[179],mul_res1[4579]);
multi_7x28 multi_7x28_mod_4580(clk,rst,matrix_A[4580],matrix_B[180],mul_res1[4580]);
multi_7x28 multi_7x28_mod_4581(clk,rst,matrix_A[4581],matrix_B[181],mul_res1[4581]);
multi_7x28 multi_7x28_mod_4582(clk,rst,matrix_A[4582],matrix_B[182],mul_res1[4582]);
multi_7x28 multi_7x28_mod_4583(clk,rst,matrix_A[4583],matrix_B[183],mul_res1[4583]);
multi_7x28 multi_7x28_mod_4584(clk,rst,matrix_A[4584],matrix_B[184],mul_res1[4584]);
multi_7x28 multi_7x28_mod_4585(clk,rst,matrix_A[4585],matrix_B[185],mul_res1[4585]);
multi_7x28 multi_7x28_mod_4586(clk,rst,matrix_A[4586],matrix_B[186],mul_res1[4586]);
multi_7x28 multi_7x28_mod_4587(clk,rst,matrix_A[4587],matrix_B[187],mul_res1[4587]);
multi_7x28 multi_7x28_mod_4588(clk,rst,matrix_A[4588],matrix_B[188],mul_res1[4588]);
multi_7x28 multi_7x28_mod_4589(clk,rst,matrix_A[4589],matrix_B[189],mul_res1[4589]);
multi_7x28 multi_7x28_mod_4590(clk,rst,matrix_A[4590],matrix_B[190],mul_res1[4590]);
multi_7x28 multi_7x28_mod_4591(clk,rst,matrix_A[4591],matrix_B[191],mul_res1[4591]);
multi_7x28 multi_7x28_mod_4592(clk,rst,matrix_A[4592],matrix_B[192],mul_res1[4592]);
multi_7x28 multi_7x28_mod_4593(clk,rst,matrix_A[4593],matrix_B[193],mul_res1[4593]);
multi_7x28 multi_7x28_mod_4594(clk,rst,matrix_A[4594],matrix_B[194],mul_res1[4594]);
multi_7x28 multi_7x28_mod_4595(clk,rst,matrix_A[4595],matrix_B[195],mul_res1[4595]);
multi_7x28 multi_7x28_mod_4596(clk,rst,matrix_A[4596],matrix_B[196],mul_res1[4596]);
multi_7x28 multi_7x28_mod_4597(clk,rst,matrix_A[4597],matrix_B[197],mul_res1[4597]);
multi_7x28 multi_7x28_mod_4598(clk,rst,matrix_A[4598],matrix_B[198],mul_res1[4598]);
multi_7x28 multi_7x28_mod_4599(clk,rst,matrix_A[4599],matrix_B[199],mul_res1[4599]);
multi_7x28 multi_7x28_mod_4600(clk,rst,matrix_A[4600],matrix_B[0],mul_res1[4600]);
multi_7x28 multi_7x28_mod_4601(clk,rst,matrix_A[4601],matrix_B[1],mul_res1[4601]);
multi_7x28 multi_7x28_mod_4602(clk,rst,matrix_A[4602],matrix_B[2],mul_res1[4602]);
multi_7x28 multi_7x28_mod_4603(clk,rst,matrix_A[4603],matrix_B[3],mul_res1[4603]);
multi_7x28 multi_7x28_mod_4604(clk,rst,matrix_A[4604],matrix_B[4],mul_res1[4604]);
multi_7x28 multi_7x28_mod_4605(clk,rst,matrix_A[4605],matrix_B[5],mul_res1[4605]);
multi_7x28 multi_7x28_mod_4606(clk,rst,matrix_A[4606],matrix_B[6],mul_res1[4606]);
multi_7x28 multi_7x28_mod_4607(clk,rst,matrix_A[4607],matrix_B[7],mul_res1[4607]);
multi_7x28 multi_7x28_mod_4608(clk,rst,matrix_A[4608],matrix_B[8],mul_res1[4608]);
multi_7x28 multi_7x28_mod_4609(clk,rst,matrix_A[4609],matrix_B[9],mul_res1[4609]);
multi_7x28 multi_7x28_mod_4610(clk,rst,matrix_A[4610],matrix_B[10],mul_res1[4610]);
multi_7x28 multi_7x28_mod_4611(clk,rst,matrix_A[4611],matrix_B[11],mul_res1[4611]);
multi_7x28 multi_7x28_mod_4612(clk,rst,matrix_A[4612],matrix_B[12],mul_res1[4612]);
multi_7x28 multi_7x28_mod_4613(clk,rst,matrix_A[4613],matrix_B[13],mul_res1[4613]);
multi_7x28 multi_7x28_mod_4614(clk,rst,matrix_A[4614],matrix_B[14],mul_res1[4614]);
multi_7x28 multi_7x28_mod_4615(clk,rst,matrix_A[4615],matrix_B[15],mul_res1[4615]);
multi_7x28 multi_7x28_mod_4616(clk,rst,matrix_A[4616],matrix_B[16],mul_res1[4616]);
multi_7x28 multi_7x28_mod_4617(clk,rst,matrix_A[4617],matrix_B[17],mul_res1[4617]);
multi_7x28 multi_7x28_mod_4618(clk,rst,matrix_A[4618],matrix_B[18],mul_res1[4618]);
multi_7x28 multi_7x28_mod_4619(clk,rst,matrix_A[4619],matrix_B[19],mul_res1[4619]);
multi_7x28 multi_7x28_mod_4620(clk,rst,matrix_A[4620],matrix_B[20],mul_res1[4620]);
multi_7x28 multi_7x28_mod_4621(clk,rst,matrix_A[4621],matrix_B[21],mul_res1[4621]);
multi_7x28 multi_7x28_mod_4622(clk,rst,matrix_A[4622],matrix_B[22],mul_res1[4622]);
multi_7x28 multi_7x28_mod_4623(clk,rst,matrix_A[4623],matrix_B[23],mul_res1[4623]);
multi_7x28 multi_7x28_mod_4624(clk,rst,matrix_A[4624],matrix_B[24],mul_res1[4624]);
multi_7x28 multi_7x28_mod_4625(clk,rst,matrix_A[4625],matrix_B[25],mul_res1[4625]);
multi_7x28 multi_7x28_mod_4626(clk,rst,matrix_A[4626],matrix_B[26],mul_res1[4626]);
multi_7x28 multi_7x28_mod_4627(clk,rst,matrix_A[4627],matrix_B[27],mul_res1[4627]);
multi_7x28 multi_7x28_mod_4628(clk,rst,matrix_A[4628],matrix_B[28],mul_res1[4628]);
multi_7x28 multi_7x28_mod_4629(clk,rst,matrix_A[4629],matrix_B[29],mul_res1[4629]);
multi_7x28 multi_7x28_mod_4630(clk,rst,matrix_A[4630],matrix_B[30],mul_res1[4630]);
multi_7x28 multi_7x28_mod_4631(clk,rst,matrix_A[4631],matrix_B[31],mul_res1[4631]);
multi_7x28 multi_7x28_mod_4632(clk,rst,matrix_A[4632],matrix_B[32],mul_res1[4632]);
multi_7x28 multi_7x28_mod_4633(clk,rst,matrix_A[4633],matrix_B[33],mul_res1[4633]);
multi_7x28 multi_7x28_mod_4634(clk,rst,matrix_A[4634],matrix_B[34],mul_res1[4634]);
multi_7x28 multi_7x28_mod_4635(clk,rst,matrix_A[4635],matrix_B[35],mul_res1[4635]);
multi_7x28 multi_7x28_mod_4636(clk,rst,matrix_A[4636],matrix_B[36],mul_res1[4636]);
multi_7x28 multi_7x28_mod_4637(clk,rst,matrix_A[4637],matrix_B[37],mul_res1[4637]);
multi_7x28 multi_7x28_mod_4638(clk,rst,matrix_A[4638],matrix_B[38],mul_res1[4638]);
multi_7x28 multi_7x28_mod_4639(clk,rst,matrix_A[4639],matrix_B[39],mul_res1[4639]);
multi_7x28 multi_7x28_mod_4640(clk,rst,matrix_A[4640],matrix_B[40],mul_res1[4640]);
multi_7x28 multi_7x28_mod_4641(clk,rst,matrix_A[4641],matrix_B[41],mul_res1[4641]);
multi_7x28 multi_7x28_mod_4642(clk,rst,matrix_A[4642],matrix_B[42],mul_res1[4642]);
multi_7x28 multi_7x28_mod_4643(clk,rst,matrix_A[4643],matrix_B[43],mul_res1[4643]);
multi_7x28 multi_7x28_mod_4644(clk,rst,matrix_A[4644],matrix_B[44],mul_res1[4644]);
multi_7x28 multi_7x28_mod_4645(clk,rst,matrix_A[4645],matrix_B[45],mul_res1[4645]);
multi_7x28 multi_7x28_mod_4646(clk,rst,matrix_A[4646],matrix_B[46],mul_res1[4646]);
multi_7x28 multi_7x28_mod_4647(clk,rst,matrix_A[4647],matrix_B[47],mul_res1[4647]);
multi_7x28 multi_7x28_mod_4648(clk,rst,matrix_A[4648],matrix_B[48],mul_res1[4648]);
multi_7x28 multi_7x28_mod_4649(clk,rst,matrix_A[4649],matrix_B[49],mul_res1[4649]);
multi_7x28 multi_7x28_mod_4650(clk,rst,matrix_A[4650],matrix_B[50],mul_res1[4650]);
multi_7x28 multi_7x28_mod_4651(clk,rst,matrix_A[4651],matrix_B[51],mul_res1[4651]);
multi_7x28 multi_7x28_mod_4652(clk,rst,matrix_A[4652],matrix_B[52],mul_res1[4652]);
multi_7x28 multi_7x28_mod_4653(clk,rst,matrix_A[4653],matrix_B[53],mul_res1[4653]);
multi_7x28 multi_7x28_mod_4654(clk,rst,matrix_A[4654],matrix_B[54],mul_res1[4654]);
multi_7x28 multi_7x28_mod_4655(clk,rst,matrix_A[4655],matrix_B[55],mul_res1[4655]);
multi_7x28 multi_7x28_mod_4656(clk,rst,matrix_A[4656],matrix_B[56],mul_res1[4656]);
multi_7x28 multi_7x28_mod_4657(clk,rst,matrix_A[4657],matrix_B[57],mul_res1[4657]);
multi_7x28 multi_7x28_mod_4658(clk,rst,matrix_A[4658],matrix_B[58],mul_res1[4658]);
multi_7x28 multi_7x28_mod_4659(clk,rst,matrix_A[4659],matrix_B[59],mul_res1[4659]);
multi_7x28 multi_7x28_mod_4660(clk,rst,matrix_A[4660],matrix_B[60],mul_res1[4660]);
multi_7x28 multi_7x28_mod_4661(clk,rst,matrix_A[4661],matrix_B[61],mul_res1[4661]);
multi_7x28 multi_7x28_mod_4662(clk,rst,matrix_A[4662],matrix_B[62],mul_res1[4662]);
multi_7x28 multi_7x28_mod_4663(clk,rst,matrix_A[4663],matrix_B[63],mul_res1[4663]);
multi_7x28 multi_7x28_mod_4664(clk,rst,matrix_A[4664],matrix_B[64],mul_res1[4664]);
multi_7x28 multi_7x28_mod_4665(clk,rst,matrix_A[4665],matrix_B[65],mul_res1[4665]);
multi_7x28 multi_7x28_mod_4666(clk,rst,matrix_A[4666],matrix_B[66],mul_res1[4666]);
multi_7x28 multi_7x28_mod_4667(clk,rst,matrix_A[4667],matrix_B[67],mul_res1[4667]);
multi_7x28 multi_7x28_mod_4668(clk,rst,matrix_A[4668],matrix_B[68],mul_res1[4668]);
multi_7x28 multi_7x28_mod_4669(clk,rst,matrix_A[4669],matrix_B[69],mul_res1[4669]);
multi_7x28 multi_7x28_mod_4670(clk,rst,matrix_A[4670],matrix_B[70],mul_res1[4670]);
multi_7x28 multi_7x28_mod_4671(clk,rst,matrix_A[4671],matrix_B[71],mul_res1[4671]);
multi_7x28 multi_7x28_mod_4672(clk,rst,matrix_A[4672],matrix_B[72],mul_res1[4672]);
multi_7x28 multi_7x28_mod_4673(clk,rst,matrix_A[4673],matrix_B[73],mul_res1[4673]);
multi_7x28 multi_7x28_mod_4674(clk,rst,matrix_A[4674],matrix_B[74],mul_res1[4674]);
multi_7x28 multi_7x28_mod_4675(clk,rst,matrix_A[4675],matrix_B[75],mul_res1[4675]);
multi_7x28 multi_7x28_mod_4676(clk,rst,matrix_A[4676],matrix_B[76],mul_res1[4676]);
multi_7x28 multi_7x28_mod_4677(clk,rst,matrix_A[4677],matrix_B[77],mul_res1[4677]);
multi_7x28 multi_7x28_mod_4678(clk,rst,matrix_A[4678],matrix_B[78],mul_res1[4678]);
multi_7x28 multi_7x28_mod_4679(clk,rst,matrix_A[4679],matrix_B[79],mul_res1[4679]);
multi_7x28 multi_7x28_mod_4680(clk,rst,matrix_A[4680],matrix_B[80],mul_res1[4680]);
multi_7x28 multi_7x28_mod_4681(clk,rst,matrix_A[4681],matrix_B[81],mul_res1[4681]);
multi_7x28 multi_7x28_mod_4682(clk,rst,matrix_A[4682],matrix_B[82],mul_res1[4682]);
multi_7x28 multi_7x28_mod_4683(clk,rst,matrix_A[4683],matrix_B[83],mul_res1[4683]);
multi_7x28 multi_7x28_mod_4684(clk,rst,matrix_A[4684],matrix_B[84],mul_res1[4684]);
multi_7x28 multi_7x28_mod_4685(clk,rst,matrix_A[4685],matrix_B[85],mul_res1[4685]);
multi_7x28 multi_7x28_mod_4686(clk,rst,matrix_A[4686],matrix_B[86],mul_res1[4686]);
multi_7x28 multi_7x28_mod_4687(clk,rst,matrix_A[4687],matrix_B[87],mul_res1[4687]);
multi_7x28 multi_7x28_mod_4688(clk,rst,matrix_A[4688],matrix_B[88],mul_res1[4688]);
multi_7x28 multi_7x28_mod_4689(clk,rst,matrix_A[4689],matrix_B[89],mul_res1[4689]);
multi_7x28 multi_7x28_mod_4690(clk,rst,matrix_A[4690],matrix_B[90],mul_res1[4690]);
multi_7x28 multi_7x28_mod_4691(clk,rst,matrix_A[4691],matrix_B[91],mul_res1[4691]);
multi_7x28 multi_7x28_mod_4692(clk,rst,matrix_A[4692],matrix_B[92],mul_res1[4692]);
multi_7x28 multi_7x28_mod_4693(clk,rst,matrix_A[4693],matrix_B[93],mul_res1[4693]);
multi_7x28 multi_7x28_mod_4694(clk,rst,matrix_A[4694],matrix_B[94],mul_res1[4694]);
multi_7x28 multi_7x28_mod_4695(clk,rst,matrix_A[4695],matrix_B[95],mul_res1[4695]);
multi_7x28 multi_7x28_mod_4696(clk,rst,matrix_A[4696],matrix_B[96],mul_res1[4696]);
multi_7x28 multi_7x28_mod_4697(clk,rst,matrix_A[4697],matrix_B[97],mul_res1[4697]);
multi_7x28 multi_7x28_mod_4698(clk,rst,matrix_A[4698],matrix_B[98],mul_res1[4698]);
multi_7x28 multi_7x28_mod_4699(clk,rst,matrix_A[4699],matrix_B[99],mul_res1[4699]);
multi_7x28 multi_7x28_mod_4700(clk,rst,matrix_A[4700],matrix_B[100],mul_res1[4700]);
multi_7x28 multi_7x28_mod_4701(clk,rst,matrix_A[4701],matrix_B[101],mul_res1[4701]);
multi_7x28 multi_7x28_mod_4702(clk,rst,matrix_A[4702],matrix_B[102],mul_res1[4702]);
multi_7x28 multi_7x28_mod_4703(clk,rst,matrix_A[4703],matrix_B[103],mul_res1[4703]);
multi_7x28 multi_7x28_mod_4704(clk,rst,matrix_A[4704],matrix_B[104],mul_res1[4704]);
multi_7x28 multi_7x28_mod_4705(clk,rst,matrix_A[4705],matrix_B[105],mul_res1[4705]);
multi_7x28 multi_7x28_mod_4706(clk,rst,matrix_A[4706],matrix_B[106],mul_res1[4706]);
multi_7x28 multi_7x28_mod_4707(clk,rst,matrix_A[4707],matrix_B[107],mul_res1[4707]);
multi_7x28 multi_7x28_mod_4708(clk,rst,matrix_A[4708],matrix_B[108],mul_res1[4708]);
multi_7x28 multi_7x28_mod_4709(clk,rst,matrix_A[4709],matrix_B[109],mul_res1[4709]);
multi_7x28 multi_7x28_mod_4710(clk,rst,matrix_A[4710],matrix_B[110],mul_res1[4710]);
multi_7x28 multi_7x28_mod_4711(clk,rst,matrix_A[4711],matrix_B[111],mul_res1[4711]);
multi_7x28 multi_7x28_mod_4712(clk,rst,matrix_A[4712],matrix_B[112],mul_res1[4712]);
multi_7x28 multi_7x28_mod_4713(clk,rst,matrix_A[4713],matrix_B[113],mul_res1[4713]);
multi_7x28 multi_7x28_mod_4714(clk,rst,matrix_A[4714],matrix_B[114],mul_res1[4714]);
multi_7x28 multi_7x28_mod_4715(clk,rst,matrix_A[4715],matrix_B[115],mul_res1[4715]);
multi_7x28 multi_7x28_mod_4716(clk,rst,matrix_A[4716],matrix_B[116],mul_res1[4716]);
multi_7x28 multi_7x28_mod_4717(clk,rst,matrix_A[4717],matrix_B[117],mul_res1[4717]);
multi_7x28 multi_7x28_mod_4718(clk,rst,matrix_A[4718],matrix_B[118],mul_res1[4718]);
multi_7x28 multi_7x28_mod_4719(clk,rst,matrix_A[4719],matrix_B[119],mul_res1[4719]);
multi_7x28 multi_7x28_mod_4720(clk,rst,matrix_A[4720],matrix_B[120],mul_res1[4720]);
multi_7x28 multi_7x28_mod_4721(clk,rst,matrix_A[4721],matrix_B[121],mul_res1[4721]);
multi_7x28 multi_7x28_mod_4722(clk,rst,matrix_A[4722],matrix_B[122],mul_res1[4722]);
multi_7x28 multi_7x28_mod_4723(clk,rst,matrix_A[4723],matrix_B[123],mul_res1[4723]);
multi_7x28 multi_7x28_mod_4724(clk,rst,matrix_A[4724],matrix_B[124],mul_res1[4724]);
multi_7x28 multi_7x28_mod_4725(clk,rst,matrix_A[4725],matrix_B[125],mul_res1[4725]);
multi_7x28 multi_7x28_mod_4726(clk,rst,matrix_A[4726],matrix_B[126],mul_res1[4726]);
multi_7x28 multi_7x28_mod_4727(clk,rst,matrix_A[4727],matrix_B[127],mul_res1[4727]);
multi_7x28 multi_7x28_mod_4728(clk,rst,matrix_A[4728],matrix_B[128],mul_res1[4728]);
multi_7x28 multi_7x28_mod_4729(clk,rst,matrix_A[4729],matrix_B[129],mul_res1[4729]);
multi_7x28 multi_7x28_mod_4730(clk,rst,matrix_A[4730],matrix_B[130],mul_res1[4730]);
multi_7x28 multi_7x28_mod_4731(clk,rst,matrix_A[4731],matrix_B[131],mul_res1[4731]);
multi_7x28 multi_7x28_mod_4732(clk,rst,matrix_A[4732],matrix_B[132],mul_res1[4732]);
multi_7x28 multi_7x28_mod_4733(clk,rst,matrix_A[4733],matrix_B[133],mul_res1[4733]);
multi_7x28 multi_7x28_mod_4734(clk,rst,matrix_A[4734],matrix_B[134],mul_res1[4734]);
multi_7x28 multi_7x28_mod_4735(clk,rst,matrix_A[4735],matrix_B[135],mul_res1[4735]);
multi_7x28 multi_7x28_mod_4736(clk,rst,matrix_A[4736],matrix_B[136],mul_res1[4736]);
multi_7x28 multi_7x28_mod_4737(clk,rst,matrix_A[4737],matrix_B[137],mul_res1[4737]);
multi_7x28 multi_7x28_mod_4738(clk,rst,matrix_A[4738],matrix_B[138],mul_res1[4738]);
multi_7x28 multi_7x28_mod_4739(clk,rst,matrix_A[4739],matrix_B[139],mul_res1[4739]);
multi_7x28 multi_7x28_mod_4740(clk,rst,matrix_A[4740],matrix_B[140],mul_res1[4740]);
multi_7x28 multi_7x28_mod_4741(clk,rst,matrix_A[4741],matrix_B[141],mul_res1[4741]);
multi_7x28 multi_7x28_mod_4742(clk,rst,matrix_A[4742],matrix_B[142],mul_res1[4742]);
multi_7x28 multi_7x28_mod_4743(clk,rst,matrix_A[4743],matrix_B[143],mul_res1[4743]);
multi_7x28 multi_7x28_mod_4744(clk,rst,matrix_A[4744],matrix_B[144],mul_res1[4744]);
multi_7x28 multi_7x28_mod_4745(clk,rst,matrix_A[4745],matrix_B[145],mul_res1[4745]);
multi_7x28 multi_7x28_mod_4746(clk,rst,matrix_A[4746],matrix_B[146],mul_res1[4746]);
multi_7x28 multi_7x28_mod_4747(clk,rst,matrix_A[4747],matrix_B[147],mul_res1[4747]);
multi_7x28 multi_7x28_mod_4748(clk,rst,matrix_A[4748],matrix_B[148],mul_res1[4748]);
multi_7x28 multi_7x28_mod_4749(clk,rst,matrix_A[4749],matrix_B[149],mul_res1[4749]);
multi_7x28 multi_7x28_mod_4750(clk,rst,matrix_A[4750],matrix_B[150],mul_res1[4750]);
multi_7x28 multi_7x28_mod_4751(clk,rst,matrix_A[4751],matrix_B[151],mul_res1[4751]);
multi_7x28 multi_7x28_mod_4752(clk,rst,matrix_A[4752],matrix_B[152],mul_res1[4752]);
multi_7x28 multi_7x28_mod_4753(clk,rst,matrix_A[4753],matrix_B[153],mul_res1[4753]);
multi_7x28 multi_7x28_mod_4754(clk,rst,matrix_A[4754],matrix_B[154],mul_res1[4754]);
multi_7x28 multi_7x28_mod_4755(clk,rst,matrix_A[4755],matrix_B[155],mul_res1[4755]);
multi_7x28 multi_7x28_mod_4756(clk,rst,matrix_A[4756],matrix_B[156],mul_res1[4756]);
multi_7x28 multi_7x28_mod_4757(clk,rst,matrix_A[4757],matrix_B[157],mul_res1[4757]);
multi_7x28 multi_7x28_mod_4758(clk,rst,matrix_A[4758],matrix_B[158],mul_res1[4758]);
multi_7x28 multi_7x28_mod_4759(clk,rst,matrix_A[4759],matrix_B[159],mul_res1[4759]);
multi_7x28 multi_7x28_mod_4760(clk,rst,matrix_A[4760],matrix_B[160],mul_res1[4760]);
multi_7x28 multi_7x28_mod_4761(clk,rst,matrix_A[4761],matrix_B[161],mul_res1[4761]);
multi_7x28 multi_7x28_mod_4762(clk,rst,matrix_A[4762],matrix_B[162],mul_res1[4762]);
multi_7x28 multi_7x28_mod_4763(clk,rst,matrix_A[4763],matrix_B[163],mul_res1[4763]);
multi_7x28 multi_7x28_mod_4764(clk,rst,matrix_A[4764],matrix_B[164],mul_res1[4764]);
multi_7x28 multi_7x28_mod_4765(clk,rst,matrix_A[4765],matrix_B[165],mul_res1[4765]);
multi_7x28 multi_7x28_mod_4766(clk,rst,matrix_A[4766],matrix_B[166],mul_res1[4766]);
multi_7x28 multi_7x28_mod_4767(clk,rst,matrix_A[4767],matrix_B[167],mul_res1[4767]);
multi_7x28 multi_7x28_mod_4768(clk,rst,matrix_A[4768],matrix_B[168],mul_res1[4768]);
multi_7x28 multi_7x28_mod_4769(clk,rst,matrix_A[4769],matrix_B[169],mul_res1[4769]);
multi_7x28 multi_7x28_mod_4770(clk,rst,matrix_A[4770],matrix_B[170],mul_res1[4770]);
multi_7x28 multi_7x28_mod_4771(clk,rst,matrix_A[4771],matrix_B[171],mul_res1[4771]);
multi_7x28 multi_7x28_mod_4772(clk,rst,matrix_A[4772],matrix_B[172],mul_res1[4772]);
multi_7x28 multi_7x28_mod_4773(clk,rst,matrix_A[4773],matrix_B[173],mul_res1[4773]);
multi_7x28 multi_7x28_mod_4774(clk,rst,matrix_A[4774],matrix_B[174],mul_res1[4774]);
multi_7x28 multi_7x28_mod_4775(clk,rst,matrix_A[4775],matrix_B[175],mul_res1[4775]);
multi_7x28 multi_7x28_mod_4776(clk,rst,matrix_A[4776],matrix_B[176],mul_res1[4776]);
multi_7x28 multi_7x28_mod_4777(clk,rst,matrix_A[4777],matrix_B[177],mul_res1[4777]);
multi_7x28 multi_7x28_mod_4778(clk,rst,matrix_A[4778],matrix_B[178],mul_res1[4778]);
multi_7x28 multi_7x28_mod_4779(clk,rst,matrix_A[4779],matrix_B[179],mul_res1[4779]);
multi_7x28 multi_7x28_mod_4780(clk,rst,matrix_A[4780],matrix_B[180],mul_res1[4780]);
multi_7x28 multi_7x28_mod_4781(clk,rst,matrix_A[4781],matrix_B[181],mul_res1[4781]);
multi_7x28 multi_7x28_mod_4782(clk,rst,matrix_A[4782],matrix_B[182],mul_res1[4782]);
multi_7x28 multi_7x28_mod_4783(clk,rst,matrix_A[4783],matrix_B[183],mul_res1[4783]);
multi_7x28 multi_7x28_mod_4784(clk,rst,matrix_A[4784],matrix_B[184],mul_res1[4784]);
multi_7x28 multi_7x28_mod_4785(clk,rst,matrix_A[4785],matrix_B[185],mul_res1[4785]);
multi_7x28 multi_7x28_mod_4786(clk,rst,matrix_A[4786],matrix_B[186],mul_res1[4786]);
multi_7x28 multi_7x28_mod_4787(clk,rst,matrix_A[4787],matrix_B[187],mul_res1[4787]);
multi_7x28 multi_7x28_mod_4788(clk,rst,matrix_A[4788],matrix_B[188],mul_res1[4788]);
multi_7x28 multi_7x28_mod_4789(clk,rst,matrix_A[4789],matrix_B[189],mul_res1[4789]);
multi_7x28 multi_7x28_mod_4790(clk,rst,matrix_A[4790],matrix_B[190],mul_res1[4790]);
multi_7x28 multi_7x28_mod_4791(clk,rst,matrix_A[4791],matrix_B[191],mul_res1[4791]);
multi_7x28 multi_7x28_mod_4792(clk,rst,matrix_A[4792],matrix_B[192],mul_res1[4792]);
multi_7x28 multi_7x28_mod_4793(clk,rst,matrix_A[4793],matrix_B[193],mul_res1[4793]);
multi_7x28 multi_7x28_mod_4794(clk,rst,matrix_A[4794],matrix_B[194],mul_res1[4794]);
multi_7x28 multi_7x28_mod_4795(clk,rst,matrix_A[4795],matrix_B[195],mul_res1[4795]);
multi_7x28 multi_7x28_mod_4796(clk,rst,matrix_A[4796],matrix_B[196],mul_res1[4796]);
multi_7x28 multi_7x28_mod_4797(clk,rst,matrix_A[4797],matrix_B[197],mul_res1[4797]);
multi_7x28 multi_7x28_mod_4798(clk,rst,matrix_A[4798],matrix_B[198],mul_res1[4798]);
multi_7x28 multi_7x28_mod_4799(clk,rst,matrix_A[4799],matrix_B[199],mul_res1[4799]);
multi_7x28 multi_7x28_mod_4800(clk,rst,matrix_A[4800],matrix_B[0],mul_res1[4800]);
multi_7x28 multi_7x28_mod_4801(clk,rst,matrix_A[4801],matrix_B[1],mul_res1[4801]);
multi_7x28 multi_7x28_mod_4802(clk,rst,matrix_A[4802],matrix_B[2],mul_res1[4802]);
multi_7x28 multi_7x28_mod_4803(clk,rst,matrix_A[4803],matrix_B[3],mul_res1[4803]);
multi_7x28 multi_7x28_mod_4804(clk,rst,matrix_A[4804],matrix_B[4],mul_res1[4804]);
multi_7x28 multi_7x28_mod_4805(clk,rst,matrix_A[4805],matrix_B[5],mul_res1[4805]);
multi_7x28 multi_7x28_mod_4806(clk,rst,matrix_A[4806],matrix_B[6],mul_res1[4806]);
multi_7x28 multi_7x28_mod_4807(clk,rst,matrix_A[4807],matrix_B[7],mul_res1[4807]);
multi_7x28 multi_7x28_mod_4808(clk,rst,matrix_A[4808],matrix_B[8],mul_res1[4808]);
multi_7x28 multi_7x28_mod_4809(clk,rst,matrix_A[4809],matrix_B[9],mul_res1[4809]);
multi_7x28 multi_7x28_mod_4810(clk,rst,matrix_A[4810],matrix_B[10],mul_res1[4810]);
multi_7x28 multi_7x28_mod_4811(clk,rst,matrix_A[4811],matrix_B[11],mul_res1[4811]);
multi_7x28 multi_7x28_mod_4812(clk,rst,matrix_A[4812],matrix_B[12],mul_res1[4812]);
multi_7x28 multi_7x28_mod_4813(clk,rst,matrix_A[4813],matrix_B[13],mul_res1[4813]);
multi_7x28 multi_7x28_mod_4814(clk,rst,matrix_A[4814],matrix_B[14],mul_res1[4814]);
multi_7x28 multi_7x28_mod_4815(clk,rst,matrix_A[4815],matrix_B[15],mul_res1[4815]);
multi_7x28 multi_7x28_mod_4816(clk,rst,matrix_A[4816],matrix_B[16],mul_res1[4816]);
multi_7x28 multi_7x28_mod_4817(clk,rst,matrix_A[4817],matrix_B[17],mul_res1[4817]);
multi_7x28 multi_7x28_mod_4818(clk,rst,matrix_A[4818],matrix_B[18],mul_res1[4818]);
multi_7x28 multi_7x28_mod_4819(clk,rst,matrix_A[4819],matrix_B[19],mul_res1[4819]);
multi_7x28 multi_7x28_mod_4820(clk,rst,matrix_A[4820],matrix_B[20],mul_res1[4820]);
multi_7x28 multi_7x28_mod_4821(clk,rst,matrix_A[4821],matrix_B[21],mul_res1[4821]);
multi_7x28 multi_7x28_mod_4822(clk,rst,matrix_A[4822],matrix_B[22],mul_res1[4822]);
multi_7x28 multi_7x28_mod_4823(clk,rst,matrix_A[4823],matrix_B[23],mul_res1[4823]);
multi_7x28 multi_7x28_mod_4824(clk,rst,matrix_A[4824],matrix_B[24],mul_res1[4824]);
multi_7x28 multi_7x28_mod_4825(clk,rst,matrix_A[4825],matrix_B[25],mul_res1[4825]);
multi_7x28 multi_7x28_mod_4826(clk,rst,matrix_A[4826],matrix_B[26],mul_res1[4826]);
multi_7x28 multi_7x28_mod_4827(clk,rst,matrix_A[4827],matrix_B[27],mul_res1[4827]);
multi_7x28 multi_7x28_mod_4828(clk,rst,matrix_A[4828],matrix_B[28],mul_res1[4828]);
multi_7x28 multi_7x28_mod_4829(clk,rst,matrix_A[4829],matrix_B[29],mul_res1[4829]);
multi_7x28 multi_7x28_mod_4830(clk,rst,matrix_A[4830],matrix_B[30],mul_res1[4830]);
multi_7x28 multi_7x28_mod_4831(clk,rst,matrix_A[4831],matrix_B[31],mul_res1[4831]);
multi_7x28 multi_7x28_mod_4832(clk,rst,matrix_A[4832],matrix_B[32],mul_res1[4832]);
multi_7x28 multi_7x28_mod_4833(clk,rst,matrix_A[4833],matrix_B[33],mul_res1[4833]);
multi_7x28 multi_7x28_mod_4834(clk,rst,matrix_A[4834],matrix_B[34],mul_res1[4834]);
multi_7x28 multi_7x28_mod_4835(clk,rst,matrix_A[4835],matrix_B[35],mul_res1[4835]);
multi_7x28 multi_7x28_mod_4836(clk,rst,matrix_A[4836],matrix_B[36],mul_res1[4836]);
multi_7x28 multi_7x28_mod_4837(clk,rst,matrix_A[4837],matrix_B[37],mul_res1[4837]);
multi_7x28 multi_7x28_mod_4838(clk,rst,matrix_A[4838],matrix_B[38],mul_res1[4838]);
multi_7x28 multi_7x28_mod_4839(clk,rst,matrix_A[4839],matrix_B[39],mul_res1[4839]);
multi_7x28 multi_7x28_mod_4840(clk,rst,matrix_A[4840],matrix_B[40],mul_res1[4840]);
multi_7x28 multi_7x28_mod_4841(clk,rst,matrix_A[4841],matrix_B[41],mul_res1[4841]);
multi_7x28 multi_7x28_mod_4842(clk,rst,matrix_A[4842],matrix_B[42],mul_res1[4842]);
multi_7x28 multi_7x28_mod_4843(clk,rst,matrix_A[4843],matrix_B[43],mul_res1[4843]);
multi_7x28 multi_7x28_mod_4844(clk,rst,matrix_A[4844],matrix_B[44],mul_res1[4844]);
multi_7x28 multi_7x28_mod_4845(clk,rst,matrix_A[4845],matrix_B[45],mul_res1[4845]);
multi_7x28 multi_7x28_mod_4846(clk,rst,matrix_A[4846],matrix_B[46],mul_res1[4846]);
multi_7x28 multi_7x28_mod_4847(clk,rst,matrix_A[4847],matrix_B[47],mul_res1[4847]);
multi_7x28 multi_7x28_mod_4848(clk,rst,matrix_A[4848],matrix_B[48],mul_res1[4848]);
multi_7x28 multi_7x28_mod_4849(clk,rst,matrix_A[4849],matrix_B[49],mul_res1[4849]);
multi_7x28 multi_7x28_mod_4850(clk,rst,matrix_A[4850],matrix_B[50],mul_res1[4850]);
multi_7x28 multi_7x28_mod_4851(clk,rst,matrix_A[4851],matrix_B[51],mul_res1[4851]);
multi_7x28 multi_7x28_mod_4852(clk,rst,matrix_A[4852],matrix_B[52],mul_res1[4852]);
multi_7x28 multi_7x28_mod_4853(clk,rst,matrix_A[4853],matrix_B[53],mul_res1[4853]);
multi_7x28 multi_7x28_mod_4854(clk,rst,matrix_A[4854],matrix_B[54],mul_res1[4854]);
multi_7x28 multi_7x28_mod_4855(clk,rst,matrix_A[4855],matrix_B[55],mul_res1[4855]);
multi_7x28 multi_7x28_mod_4856(clk,rst,matrix_A[4856],matrix_B[56],mul_res1[4856]);
multi_7x28 multi_7x28_mod_4857(clk,rst,matrix_A[4857],matrix_B[57],mul_res1[4857]);
multi_7x28 multi_7x28_mod_4858(clk,rst,matrix_A[4858],matrix_B[58],mul_res1[4858]);
multi_7x28 multi_7x28_mod_4859(clk,rst,matrix_A[4859],matrix_B[59],mul_res1[4859]);
multi_7x28 multi_7x28_mod_4860(clk,rst,matrix_A[4860],matrix_B[60],mul_res1[4860]);
multi_7x28 multi_7x28_mod_4861(clk,rst,matrix_A[4861],matrix_B[61],mul_res1[4861]);
multi_7x28 multi_7x28_mod_4862(clk,rst,matrix_A[4862],matrix_B[62],mul_res1[4862]);
multi_7x28 multi_7x28_mod_4863(clk,rst,matrix_A[4863],matrix_B[63],mul_res1[4863]);
multi_7x28 multi_7x28_mod_4864(clk,rst,matrix_A[4864],matrix_B[64],mul_res1[4864]);
multi_7x28 multi_7x28_mod_4865(clk,rst,matrix_A[4865],matrix_B[65],mul_res1[4865]);
multi_7x28 multi_7x28_mod_4866(clk,rst,matrix_A[4866],matrix_B[66],mul_res1[4866]);
multi_7x28 multi_7x28_mod_4867(clk,rst,matrix_A[4867],matrix_B[67],mul_res1[4867]);
multi_7x28 multi_7x28_mod_4868(clk,rst,matrix_A[4868],matrix_B[68],mul_res1[4868]);
multi_7x28 multi_7x28_mod_4869(clk,rst,matrix_A[4869],matrix_B[69],mul_res1[4869]);
multi_7x28 multi_7x28_mod_4870(clk,rst,matrix_A[4870],matrix_B[70],mul_res1[4870]);
multi_7x28 multi_7x28_mod_4871(clk,rst,matrix_A[4871],matrix_B[71],mul_res1[4871]);
multi_7x28 multi_7x28_mod_4872(clk,rst,matrix_A[4872],matrix_B[72],mul_res1[4872]);
multi_7x28 multi_7x28_mod_4873(clk,rst,matrix_A[4873],matrix_B[73],mul_res1[4873]);
multi_7x28 multi_7x28_mod_4874(clk,rst,matrix_A[4874],matrix_B[74],mul_res1[4874]);
multi_7x28 multi_7x28_mod_4875(clk,rst,matrix_A[4875],matrix_B[75],mul_res1[4875]);
multi_7x28 multi_7x28_mod_4876(clk,rst,matrix_A[4876],matrix_B[76],mul_res1[4876]);
multi_7x28 multi_7x28_mod_4877(clk,rst,matrix_A[4877],matrix_B[77],mul_res1[4877]);
multi_7x28 multi_7x28_mod_4878(clk,rst,matrix_A[4878],matrix_B[78],mul_res1[4878]);
multi_7x28 multi_7x28_mod_4879(clk,rst,matrix_A[4879],matrix_B[79],mul_res1[4879]);
multi_7x28 multi_7x28_mod_4880(clk,rst,matrix_A[4880],matrix_B[80],mul_res1[4880]);
multi_7x28 multi_7x28_mod_4881(clk,rst,matrix_A[4881],matrix_B[81],mul_res1[4881]);
multi_7x28 multi_7x28_mod_4882(clk,rst,matrix_A[4882],matrix_B[82],mul_res1[4882]);
multi_7x28 multi_7x28_mod_4883(clk,rst,matrix_A[4883],matrix_B[83],mul_res1[4883]);
multi_7x28 multi_7x28_mod_4884(clk,rst,matrix_A[4884],matrix_B[84],mul_res1[4884]);
multi_7x28 multi_7x28_mod_4885(clk,rst,matrix_A[4885],matrix_B[85],mul_res1[4885]);
multi_7x28 multi_7x28_mod_4886(clk,rst,matrix_A[4886],matrix_B[86],mul_res1[4886]);
multi_7x28 multi_7x28_mod_4887(clk,rst,matrix_A[4887],matrix_B[87],mul_res1[4887]);
multi_7x28 multi_7x28_mod_4888(clk,rst,matrix_A[4888],matrix_B[88],mul_res1[4888]);
multi_7x28 multi_7x28_mod_4889(clk,rst,matrix_A[4889],matrix_B[89],mul_res1[4889]);
multi_7x28 multi_7x28_mod_4890(clk,rst,matrix_A[4890],matrix_B[90],mul_res1[4890]);
multi_7x28 multi_7x28_mod_4891(clk,rst,matrix_A[4891],matrix_B[91],mul_res1[4891]);
multi_7x28 multi_7x28_mod_4892(clk,rst,matrix_A[4892],matrix_B[92],mul_res1[4892]);
multi_7x28 multi_7x28_mod_4893(clk,rst,matrix_A[4893],matrix_B[93],mul_res1[4893]);
multi_7x28 multi_7x28_mod_4894(clk,rst,matrix_A[4894],matrix_B[94],mul_res1[4894]);
multi_7x28 multi_7x28_mod_4895(clk,rst,matrix_A[4895],matrix_B[95],mul_res1[4895]);
multi_7x28 multi_7x28_mod_4896(clk,rst,matrix_A[4896],matrix_B[96],mul_res1[4896]);
multi_7x28 multi_7x28_mod_4897(clk,rst,matrix_A[4897],matrix_B[97],mul_res1[4897]);
multi_7x28 multi_7x28_mod_4898(clk,rst,matrix_A[4898],matrix_B[98],mul_res1[4898]);
multi_7x28 multi_7x28_mod_4899(clk,rst,matrix_A[4899],matrix_B[99],mul_res1[4899]);
multi_7x28 multi_7x28_mod_4900(clk,rst,matrix_A[4900],matrix_B[100],mul_res1[4900]);
multi_7x28 multi_7x28_mod_4901(clk,rst,matrix_A[4901],matrix_B[101],mul_res1[4901]);
multi_7x28 multi_7x28_mod_4902(clk,rst,matrix_A[4902],matrix_B[102],mul_res1[4902]);
multi_7x28 multi_7x28_mod_4903(clk,rst,matrix_A[4903],matrix_B[103],mul_res1[4903]);
multi_7x28 multi_7x28_mod_4904(clk,rst,matrix_A[4904],matrix_B[104],mul_res1[4904]);
multi_7x28 multi_7x28_mod_4905(clk,rst,matrix_A[4905],matrix_B[105],mul_res1[4905]);
multi_7x28 multi_7x28_mod_4906(clk,rst,matrix_A[4906],matrix_B[106],mul_res1[4906]);
multi_7x28 multi_7x28_mod_4907(clk,rst,matrix_A[4907],matrix_B[107],mul_res1[4907]);
multi_7x28 multi_7x28_mod_4908(clk,rst,matrix_A[4908],matrix_B[108],mul_res1[4908]);
multi_7x28 multi_7x28_mod_4909(clk,rst,matrix_A[4909],matrix_B[109],mul_res1[4909]);
multi_7x28 multi_7x28_mod_4910(clk,rst,matrix_A[4910],matrix_B[110],mul_res1[4910]);
multi_7x28 multi_7x28_mod_4911(clk,rst,matrix_A[4911],matrix_B[111],mul_res1[4911]);
multi_7x28 multi_7x28_mod_4912(clk,rst,matrix_A[4912],matrix_B[112],mul_res1[4912]);
multi_7x28 multi_7x28_mod_4913(clk,rst,matrix_A[4913],matrix_B[113],mul_res1[4913]);
multi_7x28 multi_7x28_mod_4914(clk,rst,matrix_A[4914],matrix_B[114],mul_res1[4914]);
multi_7x28 multi_7x28_mod_4915(clk,rst,matrix_A[4915],matrix_B[115],mul_res1[4915]);
multi_7x28 multi_7x28_mod_4916(clk,rst,matrix_A[4916],matrix_B[116],mul_res1[4916]);
multi_7x28 multi_7x28_mod_4917(clk,rst,matrix_A[4917],matrix_B[117],mul_res1[4917]);
multi_7x28 multi_7x28_mod_4918(clk,rst,matrix_A[4918],matrix_B[118],mul_res1[4918]);
multi_7x28 multi_7x28_mod_4919(clk,rst,matrix_A[4919],matrix_B[119],mul_res1[4919]);
multi_7x28 multi_7x28_mod_4920(clk,rst,matrix_A[4920],matrix_B[120],mul_res1[4920]);
multi_7x28 multi_7x28_mod_4921(clk,rst,matrix_A[4921],matrix_B[121],mul_res1[4921]);
multi_7x28 multi_7x28_mod_4922(clk,rst,matrix_A[4922],matrix_B[122],mul_res1[4922]);
multi_7x28 multi_7x28_mod_4923(clk,rst,matrix_A[4923],matrix_B[123],mul_res1[4923]);
multi_7x28 multi_7x28_mod_4924(clk,rst,matrix_A[4924],matrix_B[124],mul_res1[4924]);
multi_7x28 multi_7x28_mod_4925(clk,rst,matrix_A[4925],matrix_B[125],mul_res1[4925]);
multi_7x28 multi_7x28_mod_4926(clk,rst,matrix_A[4926],matrix_B[126],mul_res1[4926]);
multi_7x28 multi_7x28_mod_4927(clk,rst,matrix_A[4927],matrix_B[127],mul_res1[4927]);
multi_7x28 multi_7x28_mod_4928(clk,rst,matrix_A[4928],matrix_B[128],mul_res1[4928]);
multi_7x28 multi_7x28_mod_4929(clk,rst,matrix_A[4929],matrix_B[129],mul_res1[4929]);
multi_7x28 multi_7x28_mod_4930(clk,rst,matrix_A[4930],matrix_B[130],mul_res1[4930]);
multi_7x28 multi_7x28_mod_4931(clk,rst,matrix_A[4931],matrix_B[131],mul_res1[4931]);
multi_7x28 multi_7x28_mod_4932(clk,rst,matrix_A[4932],matrix_B[132],mul_res1[4932]);
multi_7x28 multi_7x28_mod_4933(clk,rst,matrix_A[4933],matrix_B[133],mul_res1[4933]);
multi_7x28 multi_7x28_mod_4934(clk,rst,matrix_A[4934],matrix_B[134],mul_res1[4934]);
multi_7x28 multi_7x28_mod_4935(clk,rst,matrix_A[4935],matrix_B[135],mul_res1[4935]);
multi_7x28 multi_7x28_mod_4936(clk,rst,matrix_A[4936],matrix_B[136],mul_res1[4936]);
multi_7x28 multi_7x28_mod_4937(clk,rst,matrix_A[4937],matrix_B[137],mul_res1[4937]);
multi_7x28 multi_7x28_mod_4938(clk,rst,matrix_A[4938],matrix_B[138],mul_res1[4938]);
multi_7x28 multi_7x28_mod_4939(clk,rst,matrix_A[4939],matrix_B[139],mul_res1[4939]);
multi_7x28 multi_7x28_mod_4940(clk,rst,matrix_A[4940],matrix_B[140],mul_res1[4940]);
multi_7x28 multi_7x28_mod_4941(clk,rst,matrix_A[4941],matrix_B[141],mul_res1[4941]);
multi_7x28 multi_7x28_mod_4942(clk,rst,matrix_A[4942],matrix_B[142],mul_res1[4942]);
multi_7x28 multi_7x28_mod_4943(clk,rst,matrix_A[4943],matrix_B[143],mul_res1[4943]);
multi_7x28 multi_7x28_mod_4944(clk,rst,matrix_A[4944],matrix_B[144],mul_res1[4944]);
multi_7x28 multi_7x28_mod_4945(clk,rst,matrix_A[4945],matrix_B[145],mul_res1[4945]);
multi_7x28 multi_7x28_mod_4946(clk,rst,matrix_A[4946],matrix_B[146],mul_res1[4946]);
multi_7x28 multi_7x28_mod_4947(clk,rst,matrix_A[4947],matrix_B[147],mul_res1[4947]);
multi_7x28 multi_7x28_mod_4948(clk,rst,matrix_A[4948],matrix_B[148],mul_res1[4948]);
multi_7x28 multi_7x28_mod_4949(clk,rst,matrix_A[4949],matrix_B[149],mul_res1[4949]);
multi_7x28 multi_7x28_mod_4950(clk,rst,matrix_A[4950],matrix_B[150],mul_res1[4950]);
multi_7x28 multi_7x28_mod_4951(clk,rst,matrix_A[4951],matrix_B[151],mul_res1[4951]);
multi_7x28 multi_7x28_mod_4952(clk,rst,matrix_A[4952],matrix_B[152],mul_res1[4952]);
multi_7x28 multi_7x28_mod_4953(clk,rst,matrix_A[4953],matrix_B[153],mul_res1[4953]);
multi_7x28 multi_7x28_mod_4954(clk,rst,matrix_A[4954],matrix_B[154],mul_res1[4954]);
multi_7x28 multi_7x28_mod_4955(clk,rst,matrix_A[4955],matrix_B[155],mul_res1[4955]);
multi_7x28 multi_7x28_mod_4956(clk,rst,matrix_A[4956],matrix_B[156],mul_res1[4956]);
multi_7x28 multi_7x28_mod_4957(clk,rst,matrix_A[4957],matrix_B[157],mul_res1[4957]);
multi_7x28 multi_7x28_mod_4958(clk,rst,matrix_A[4958],matrix_B[158],mul_res1[4958]);
multi_7x28 multi_7x28_mod_4959(clk,rst,matrix_A[4959],matrix_B[159],mul_res1[4959]);
multi_7x28 multi_7x28_mod_4960(clk,rst,matrix_A[4960],matrix_B[160],mul_res1[4960]);
multi_7x28 multi_7x28_mod_4961(clk,rst,matrix_A[4961],matrix_B[161],mul_res1[4961]);
multi_7x28 multi_7x28_mod_4962(clk,rst,matrix_A[4962],matrix_B[162],mul_res1[4962]);
multi_7x28 multi_7x28_mod_4963(clk,rst,matrix_A[4963],matrix_B[163],mul_res1[4963]);
multi_7x28 multi_7x28_mod_4964(clk,rst,matrix_A[4964],matrix_B[164],mul_res1[4964]);
multi_7x28 multi_7x28_mod_4965(clk,rst,matrix_A[4965],matrix_B[165],mul_res1[4965]);
multi_7x28 multi_7x28_mod_4966(clk,rst,matrix_A[4966],matrix_B[166],mul_res1[4966]);
multi_7x28 multi_7x28_mod_4967(clk,rst,matrix_A[4967],matrix_B[167],mul_res1[4967]);
multi_7x28 multi_7x28_mod_4968(clk,rst,matrix_A[4968],matrix_B[168],mul_res1[4968]);
multi_7x28 multi_7x28_mod_4969(clk,rst,matrix_A[4969],matrix_B[169],mul_res1[4969]);
multi_7x28 multi_7x28_mod_4970(clk,rst,matrix_A[4970],matrix_B[170],mul_res1[4970]);
multi_7x28 multi_7x28_mod_4971(clk,rst,matrix_A[4971],matrix_B[171],mul_res1[4971]);
multi_7x28 multi_7x28_mod_4972(clk,rst,matrix_A[4972],matrix_B[172],mul_res1[4972]);
multi_7x28 multi_7x28_mod_4973(clk,rst,matrix_A[4973],matrix_B[173],mul_res1[4973]);
multi_7x28 multi_7x28_mod_4974(clk,rst,matrix_A[4974],matrix_B[174],mul_res1[4974]);
multi_7x28 multi_7x28_mod_4975(clk,rst,matrix_A[4975],matrix_B[175],mul_res1[4975]);
multi_7x28 multi_7x28_mod_4976(clk,rst,matrix_A[4976],matrix_B[176],mul_res1[4976]);
multi_7x28 multi_7x28_mod_4977(clk,rst,matrix_A[4977],matrix_B[177],mul_res1[4977]);
multi_7x28 multi_7x28_mod_4978(clk,rst,matrix_A[4978],matrix_B[178],mul_res1[4978]);
multi_7x28 multi_7x28_mod_4979(clk,rst,matrix_A[4979],matrix_B[179],mul_res1[4979]);
multi_7x28 multi_7x28_mod_4980(clk,rst,matrix_A[4980],matrix_B[180],mul_res1[4980]);
multi_7x28 multi_7x28_mod_4981(clk,rst,matrix_A[4981],matrix_B[181],mul_res1[4981]);
multi_7x28 multi_7x28_mod_4982(clk,rst,matrix_A[4982],matrix_B[182],mul_res1[4982]);
multi_7x28 multi_7x28_mod_4983(clk,rst,matrix_A[4983],matrix_B[183],mul_res1[4983]);
multi_7x28 multi_7x28_mod_4984(clk,rst,matrix_A[4984],matrix_B[184],mul_res1[4984]);
multi_7x28 multi_7x28_mod_4985(clk,rst,matrix_A[4985],matrix_B[185],mul_res1[4985]);
multi_7x28 multi_7x28_mod_4986(clk,rst,matrix_A[4986],matrix_B[186],mul_res1[4986]);
multi_7x28 multi_7x28_mod_4987(clk,rst,matrix_A[4987],matrix_B[187],mul_res1[4987]);
multi_7x28 multi_7x28_mod_4988(clk,rst,matrix_A[4988],matrix_B[188],mul_res1[4988]);
multi_7x28 multi_7x28_mod_4989(clk,rst,matrix_A[4989],matrix_B[189],mul_res1[4989]);
multi_7x28 multi_7x28_mod_4990(clk,rst,matrix_A[4990],matrix_B[190],mul_res1[4990]);
multi_7x28 multi_7x28_mod_4991(clk,rst,matrix_A[4991],matrix_B[191],mul_res1[4991]);
multi_7x28 multi_7x28_mod_4992(clk,rst,matrix_A[4992],matrix_B[192],mul_res1[4992]);
multi_7x28 multi_7x28_mod_4993(clk,rst,matrix_A[4993],matrix_B[193],mul_res1[4993]);
multi_7x28 multi_7x28_mod_4994(clk,rst,matrix_A[4994],matrix_B[194],mul_res1[4994]);
multi_7x28 multi_7x28_mod_4995(clk,rst,matrix_A[4995],matrix_B[195],mul_res1[4995]);
multi_7x28 multi_7x28_mod_4996(clk,rst,matrix_A[4996],matrix_B[196],mul_res1[4996]);
multi_7x28 multi_7x28_mod_4997(clk,rst,matrix_A[4997],matrix_B[197],mul_res1[4997]);
multi_7x28 multi_7x28_mod_4998(clk,rst,matrix_A[4998],matrix_B[198],mul_res1[4998]);
multi_7x28 multi_7x28_mod_4999(clk,rst,matrix_A[4999],matrix_B[199],mul_res1[4999]);
multi_7x28 multi_7x28_mod_5000(clk,rst,matrix_A[5000],matrix_B[0],mul_res1[5000]);
multi_7x28 multi_7x28_mod_5001(clk,rst,matrix_A[5001],matrix_B[1],mul_res1[5001]);
multi_7x28 multi_7x28_mod_5002(clk,rst,matrix_A[5002],matrix_B[2],mul_res1[5002]);
multi_7x28 multi_7x28_mod_5003(clk,rst,matrix_A[5003],matrix_B[3],mul_res1[5003]);
multi_7x28 multi_7x28_mod_5004(clk,rst,matrix_A[5004],matrix_B[4],mul_res1[5004]);
multi_7x28 multi_7x28_mod_5005(clk,rst,matrix_A[5005],matrix_B[5],mul_res1[5005]);
multi_7x28 multi_7x28_mod_5006(clk,rst,matrix_A[5006],matrix_B[6],mul_res1[5006]);
multi_7x28 multi_7x28_mod_5007(clk,rst,matrix_A[5007],matrix_B[7],mul_res1[5007]);
multi_7x28 multi_7x28_mod_5008(clk,rst,matrix_A[5008],matrix_B[8],mul_res1[5008]);
multi_7x28 multi_7x28_mod_5009(clk,rst,matrix_A[5009],matrix_B[9],mul_res1[5009]);
multi_7x28 multi_7x28_mod_5010(clk,rst,matrix_A[5010],matrix_B[10],mul_res1[5010]);
multi_7x28 multi_7x28_mod_5011(clk,rst,matrix_A[5011],matrix_B[11],mul_res1[5011]);
multi_7x28 multi_7x28_mod_5012(clk,rst,matrix_A[5012],matrix_B[12],mul_res1[5012]);
multi_7x28 multi_7x28_mod_5013(clk,rst,matrix_A[5013],matrix_B[13],mul_res1[5013]);
multi_7x28 multi_7x28_mod_5014(clk,rst,matrix_A[5014],matrix_B[14],mul_res1[5014]);
multi_7x28 multi_7x28_mod_5015(clk,rst,matrix_A[5015],matrix_B[15],mul_res1[5015]);
multi_7x28 multi_7x28_mod_5016(clk,rst,matrix_A[5016],matrix_B[16],mul_res1[5016]);
multi_7x28 multi_7x28_mod_5017(clk,rst,matrix_A[5017],matrix_B[17],mul_res1[5017]);
multi_7x28 multi_7x28_mod_5018(clk,rst,matrix_A[5018],matrix_B[18],mul_res1[5018]);
multi_7x28 multi_7x28_mod_5019(clk,rst,matrix_A[5019],matrix_B[19],mul_res1[5019]);
multi_7x28 multi_7x28_mod_5020(clk,rst,matrix_A[5020],matrix_B[20],mul_res1[5020]);
multi_7x28 multi_7x28_mod_5021(clk,rst,matrix_A[5021],matrix_B[21],mul_res1[5021]);
multi_7x28 multi_7x28_mod_5022(clk,rst,matrix_A[5022],matrix_B[22],mul_res1[5022]);
multi_7x28 multi_7x28_mod_5023(clk,rst,matrix_A[5023],matrix_B[23],mul_res1[5023]);
multi_7x28 multi_7x28_mod_5024(clk,rst,matrix_A[5024],matrix_B[24],mul_res1[5024]);
multi_7x28 multi_7x28_mod_5025(clk,rst,matrix_A[5025],matrix_B[25],mul_res1[5025]);
multi_7x28 multi_7x28_mod_5026(clk,rst,matrix_A[5026],matrix_B[26],mul_res1[5026]);
multi_7x28 multi_7x28_mod_5027(clk,rst,matrix_A[5027],matrix_B[27],mul_res1[5027]);
multi_7x28 multi_7x28_mod_5028(clk,rst,matrix_A[5028],matrix_B[28],mul_res1[5028]);
multi_7x28 multi_7x28_mod_5029(clk,rst,matrix_A[5029],matrix_B[29],mul_res1[5029]);
multi_7x28 multi_7x28_mod_5030(clk,rst,matrix_A[5030],matrix_B[30],mul_res1[5030]);
multi_7x28 multi_7x28_mod_5031(clk,rst,matrix_A[5031],matrix_B[31],mul_res1[5031]);
multi_7x28 multi_7x28_mod_5032(clk,rst,matrix_A[5032],matrix_B[32],mul_res1[5032]);
multi_7x28 multi_7x28_mod_5033(clk,rst,matrix_A[5033],matrix_B[33],mul_res1[5033]);
multi_7x28 multi_7x28_mod_5034(clk,rst,matrix_A[5034],matrix_B[34],mul_res1[5034]);
multi_7x28 multi_7x28_mod_5035(clk,rst,matrix_A[5035],matrix_B[35],mul_res1[5035]);
multi_7x28 multi_7x28_mod_5036(clk,rst,matrix_A[5036],matrix_B[36],mul_res1[5036]);
multi_7x28 multi_7x28_mod_5037(clk,rst,matrix_A[5037],matrix_B[37],mul_res1[5037]);
multi_7x28 multi_7x28_mod_5038(clk,rst,matrix_A[5038],matrix_B[38],mul_res1[5038]);
multi_7x28 multi_7x28_mod_5039(clk,rst,matrix_A[5039],matrix_B[39],mul_res1[5039]);
multi_7x28 multi_7x28_mod_5040(clk,rst,matrix_A[5040],matrix_B[40],mul_res1[5040]);
multi_7x28 multi_7x28_mod_5041(clk,rst,matrix_A[5041],matrix_B[41],mul_res1[5041]);
multi_7x28 multi_7x28_mod_5042(clk,rst,matrix_A[5042],matrix_B[42],mul_res1[5042]);
multi_7x28 multi_7x28_mod_5043(clk,rst,matrix_A[5043],matrix_B[43],mul_res1[5043]);
multi_7x28 multi_7x28_mod_5044(clk,rst,matrix_A[5044],matrix_B[44],mul_res1[5044]);
multi_7x28 multi_7x28_mod_5045(clk,rst,matrix_A[5045],matrix_B[45],mul_res1[5045]);
multi_7x28 multi_7x28_mod_5046(clk,rst,matrix_A[5046],matrix_B[46],mul_res1[5046]);
multi_7x28 multi_7x28_mod_5047(clk,rst,matrix_A[5047],matrix_B[47],mul_res1[5047]);
multi_7x28 multi_7x28_mod_5048(clk,rst,matrix_A[5048],matrix_B[48],mul_res1[5048]);
multi_7x28 multi_7x28_mod_5049(clk,rst,matrix_A[5049],matrix_B[49],mul_res1[5049]);
multi_7x28 multi_7x28_mod_5050(clk,rst,matrix_A[5050],matrix_B[50],mul_res1[5050]);
multi_7x28 multi_7x28_mod_5051(clk,rst,matrix_A[5051],matrix_B[51],mul_res1[5051]);
multi_7x28 multi_7x28_mod_5052(clk,rst,matrix_A[5052],matrix_B[52],mul_res1[5052]);
multi_7x28 multi_7x28_mod_5053(clk,rst,matrix_A[5053],matrix_B[53],mul_res1[5053]);
multi_7x28 multi_7x28_mod_5054(clk,rst,matrix_A[5054],matrix_B[54],mul_res1[5054]);
multi_7x28 multi_7x28_mod_5055(clk,rst,matrix_A[5055],matrix_B[55],mul_res1[5055]);
multi_7x28 multi_7x28_mod_5056(clk,rst,matrix_A[5056],matrix_B[56],mul_res1[5056]);
multi_7x28 multi_7x28_mod_5057(clk,rst,matrix_A[5057],matrix_B[57],mul_res1[5057]);
multi_7x28 multi_7x28_mod_5058(clk,rst,matrix_A[5058],matrix_B[58],mul_res1[5058]);
multi_7x28 multi_7x28_mod_5059(clk,rst,matrix_A[5059],matrix_B[59],mul_res1[5059]);
multi_7x28 multi_7x28_mod_5060(clk,rst,matrix_A[5060],matrix_B[60],mul_res1[5060]);
multi_7x28 multi_7x28_mod_5061(clk,rst,matrix_A[5061],matrix_B[61],mul_res1[5061]);
multi_7x28 multi_7x28_mod_5062(clk,rst,matrix_A[5062],matrix_B[62],mul_res1[5062]);
multi_7x28 multi_7x28_mod_5063(clk,rst,matrix_A[5063],matrix_B[63],mul_res1[5063]);
multi_7x28 multi_7x28_mod_5064(clk,rst,matrix_A[5064],matrix_B[64],mul_res1[5064]);
multi_7x28 multi_7x28_mod_5065(clk,rst,matrix_A[5065],matrix_B[65],mul_res1[5065]);
multi_7x28 multi_7x28_mod_5066(clk,rst,matrix_A[5066],matrix_B[66],mul_res1[5066]);
multi_7x28 multi_7x28_mod_5067(clk,rst,matrix_A[5067],matrix_B[67],mul_res1[5067]);
multi_7x28 multi_7x28_mod_5068(clk,rst,matrix_A[5068],matrix_B[68],mul_res1[5068]);
multi_7x28 multi_7x28_mod_5069(clk,rst,matrix_A[5069],matrix_B[69],mul_res1[5069]);
multi_7x28 multi_7x28_mod_5070(clk,rst,matrix_A[5070],matrix_B[70],mul_res1[5070]);
multi_7x28 multi_7x28_mod_5071(clk,rst,matrix_A[5071],matrix_B[71],mul_res1[5071]);
multi_7x28 multi_7x28_mod_5072(clk,rst,matrix_A[5072],matrix_B[72],mul_res1[5072]);
multi_7x28 multi_7x28_mod_5073(clk,rst,matrix_A[5073],matrix_B[73],mul_res1[5073]);
multi_7x28 multi_7x28_mod_5074(clk,rst,matrix_A[5074],matrix_B[74],mul_res1[5074]);
multi_7x28 multi_7x28_mod_5075(clk,rst,matrix_A[5075],matrix_B[75],mul_res1[5075]);
multi_7x28 multi_7x28_mod_5076(clk,rst,matrix_A[5076],matrix_B[76],mul_res1[5076]);
multi_7x28 multi_7x28_mod_5077(clk,rst,matrix_A[5077],matrix_B[77],mul_res1[5077]);
multi_7x28 multi_7x28_mod_5078(clk,rst,matrix_A[5078],matrix_B[78],mul_res1[5078]);
multi_7x28 multi_7x28_mod_5079(clk,rst,matrix_A[5079],matrix_B[79],mul_res1[5079]);
multi_7x28 multi_7x28_mod_5080(clk,rst,matrix_A[5080],matrix_B[80],mul_res1[5080]);
multi_7x28 multi_7x28_mod_5081(clk,rst,matrix_A[5081],matrix_B[81],mul_res1[5081]);
multi_7x28 multi_7x28_mod_5082(clk,rst,matrix_A[5082],matrix_B[82],mul_res1[5082]);
multi_7x28 multi_7x28_mod_5083(clk,rst,matrix_A[5083],matrix_B[83],mul_res1[5083]);
multi_7x28 multi_7x28_mod_5084(clk,rst,matrix_A[5084],matrix_B[84],mul_res1[5084]);
multi_7x28 multi_7x28_mod_5085(clk,rst,matrix_A[5085],matrix_B[85],mul_res1[5085]);
multi_7x28 multi_7x28_mod_5086(clk,rst,matrix_A[5086],matrix_B[86],mul_res1[5086]);
multi_7x28 multi_7x28_mod_5087(clk,rst,matrix_A[5087],matrix_B[87],mul_res1[5087]);
multi_7x28 multi_7x28_mod_5088(clk,rst,matrix_A[5088],matrix_B[88],mul_res1[5088]);
multi_7x28 multi_7x28_mod_5089(clk,rst,matrix_A[5089],matrix_B[89],mul_res1[5089]);
multi_7x28 multi_7x28_mod_5090(clk,rst,matrix_A[5090],matrix_B[90],mul_res1[5090]);
multi_7x28 multi_7x28_mod_5091(clk,rst,matrix_A[5091],matrix_B[91],mul_res1[5091]);
multi_7x28 multi_7x28_mod_5092(clk,rst,matrix_A[5092],matrix_B[92],mul_res1[5092]);
multi_7x28 multi_7x28_mod_5093(clk,rst,matrix_A[5093],matrix_B[93],mul_res1[5093]);
multi_7x28 multi_7x28_mod_5094(clk,rst,matrix_A[5094],matrix_B[94],mul_res1[5094]);
multi_7x28 multi_7x28_mod_5095(clk,rst,matrix_A[5095],matrix_B[95],mul_res1[5095]);
multi_7x28 multi_7x28_mod_5096(clk,rst,matrix_A[5096],matrix_B[96],mul_res1[5096]);
multi_7x28 multi_7x28_mod_5097(clk,rst,matrix_A[5097],matrix_B[97],mul_res1[5097]);
multi_7x28 multi_7x28_mod_5098(clk,rst,matrix_A[5098],matrix_B[98],mul_res1[5098]);
multi_7x28 multi_7x28_mod_5099(clk,rst,matrix_A[5099],matrix_B[99],mul_res1[5099]);
multi_7x28 multi_7x28_mod_5100(clk,rst,matrix_A[5100],matrix_B[100],mul_res1[5100]);
multi_7x28 multi_7x28_mod_5101(clk,rst,matrix_A[5101],matrix_B[101],mul_res1[5101]);
multi_7x28 multi_7x28_mod_5102(clk,rst,matrix_A[5102],matrix_B[102],mul_res1[5102]);
multi_7x28 multi_7x28_mod_5103(clk,rst,matrix_A[5103],matrix_B[103],mul_res1[5103]);
multi_7x28 multi_7x28_mod_5104(clk,rst,matrix_A[5104],matrix_B[104],mul_res1[5104]);
multi_7x28 multi_7x28_mod_5105(clk,rst,matrix_A[5105],matrix_B[105],mul_res1[5105]);
multi_7x28 multi_7x28_mod_5106(clk,rst,matrix_A[5106],matrix_B[106],mul_res1[5106]);
multi_7x28 multi_7x28_mod_5107(clk,rst,matrix_A[5107],matrix_B[107],mul_res1[5107]);
multi_7x28 multi_7x28_mod_5108(clk,rst,matrix_A[5108],matrix_B[108],mul_res1[5108]);
multi_7x28 multi_7x28_mod_5109(clk,rst,matrix_A[5109],matrix_B[109],mul_res1[5109]);
multi_7x28 multi_7x28_mod_5110(clk,rst,matrix_A[5110],matrix_B[110],mul_res1[5110]);
multi_7x28 multi_7x28_mod_5111(clk,rst,matrix_A[5111],matrix_B[111],mul_res1[5111]);
multi_7x28 multi_7x28_mod_5112(clk,rst,matrix_A[5112],matrix_B[112],mul_res1[5112]);
multi_7x28 multi_7x28_mod_5113(clk,rst,matrix_A[5113],matrix_B[113],mul_res1[5113]);
multi_7x28 multi_7x28_mod_5114(clk,rst,matrix_A[5114],matrix_B[114],mul_res1[5114]);
multi_7x28 multi_7x28_mod_5115(clk,rst,matrix_A[5115],matrix_B[115],mul_res1[5115]);
multi_7x28 multi_7x28_mod_5116(clk,rst,matrix_A[5116],matrix_B[116],mul_res1[5116]);
multi_7x28 multi_7x28_mod_5117(clk,rst,matrix_A[5117],matrix_B[117],mul_res1[5117]);
multi_7x28 multi_7x28_mod_5118(clk,rst,matrix_A[5118],matrix_B[118],mul_res1[5118]);
multi_7x28 multi_7x28_mod_5119(clk,rst,matrix_A[5119],matrix_B[119],mul_res1[5119]);
multi_7x28 multi_7x28_mod_5120(clk,rst,matrix_A[5120],matrix_B[120],mul_res1[5120]);
multi_7x28 multi_7x28_mod_5121(clk,rst,matrix_A[5121],matrix_B[121],mul_res1[5121]);
multi_7x28 multi_7x28_mod_5122(clk,rst,matrix_A[5122],matrix_B[122],mul_res1[5122]);
multi_7x28 multi_7x28_mod_5123(clk,rst,matrix_A[5123],matrix_B[123],mul_res1[5123]);
multi_7x28 multi_7x28_mod_5124(clk,rst,matrix_A[5124],matrix_B[124],mul_res1[5124]);
multi_7x28 multi_7x28_mod_5125(clk,rst,matrix_A[5125],matrix_B[125],mul_res1[5125]);
multi_7x28 multi_7x28_mod_5126(clk,rst,matrix_A[5126],matrix_B[126],mul_res1[5126]);
multi_7x28 multi_7x28_mod_5127(clk,rst,matrix_A[5127],matrix_B[127],mul_res1[5127]);
multi_7x28 multi_7x28_mod_5128(clk,rst,matrix_A[5128],matrix_B[128],mul_res1[5128]);
multi_7x28 multi_7x28_mod_5129(clk,rst,matrix_A[5129],matrix_B[129],mul_res1[5129]);
multi_7x28 multi_7x28_mod_5130(clk,rst,matrix_A[5130],matrix_B[130],mul_res1[5130]);
multi_7x28 multi_7x28_mod_5131(clk,rst,matrix_A[5131],matrix_B[131],mul_res1[5131]);
multi_7x28 multi_7x28_mod_5132(clk,rst,matrix_A[5132],matrix_B[132],mul_res1[5132]);
multi_7x28 multi_7x28_mod_5133(clk,rst,matrix_A[5133],matrix_B[133],mul_res1[5133]);
multi_7x28 multi_7x28_mod_5134(clk,rst,matrix_A[5134],matrix_B[134],mul_res1[5134]);
multi_7x28 multi_7x28_mod_5135(clk,rst,matrix_A[5135],matrix_B[135],mul_res1[5135]);
multi_7x28 multi_7x28_mod_5136(clk,rst,matrix_A[5136],matrix_B[136],mul_res1[5136]);
multi_7x28 multi_7x28_mod_5137(clk,rst,matrix_A[5137],matrix_B[137],mul_res1[5137]);
multi_7x28 multi_7x28_mod_5138(clk,rst,matrix_A[5138],matrix_B[138],mul_res1[5138]);
multi_7x28 multi_7x28_mod_5139(clk,rst,matrix_A[5139],matrix_B[139],mul_res1[5139]);
multi_7x28 multi_7x28_mod_5140(clk,rst,matrix_A[5140],matrix_B[140],mul_res1[5140]);
multi_7x28 multi_7x28_mod_5141(clk,rst,matrix_A[5141],matrix_B[141],mul_res1[5141]);
multi_7x28 multi_7x28_mod_5142(clk,rst,matrix_A[5142],matrix_B[142],mul_res1[5142]);
multi_7x28 multi_7x28_mod_5143(clk,rst,matrix_A[5143],matrix_B[143],mul_res1[5143]);
multi_7x28 multi_7x28_mod_5144(clk,rst,matrix_A[5144],matrix_B[144],mul_res1[5144]);
multi_7x28 multi_7x28_mod_5145(clk,rst,matrix_A[5145],matrix_B[145],mul_res1[5145]);
multi_7x28 multi_7x28_mod_5146(clk,rst,matrix_A[5146],matrix_B[146],mul_res1[5146]);
multi_7x28 multi_7x28_mod_5147(clk,rst,matrix_A[5147],matrix_B[147],mul_res1[5147]);
multi_7x28 multi_7x28_mod_5148(clk,rst,matrix_A[5148],matrix_B[148],mul_res1[5148]);
multi_7x28 multi_7x28_mod_5149(clk,rst,matrix_A[5149],matrix_B[149],mul_res1[5149]);
multi_7x28 multi_7x28_mod_5150(clk,rst,matrix_A[5150],matrix_B[150],mul_res1[5150]);
multi_7x28 multi_7x28_mod_5151(clk,rst,matrix_A[5151],matrix_B[151],mul_res1[5151]);
multi_7x28 multi_7x28_mod_5152(clk,rst,matrix_A[5152],matrix_B[152],mul_res1[5152]);
multi_7x28 multi_7x28_mod_5153(clk,rst,matrix_A[5153],matrix_B[153],mul_res1[5153]);
multi_7x28 multi_7x28_mod_5154(clk,rst,matrix_A[5154],matrix_B[154],mul_res1[5154]);
multi_7x28 multi_7x28_mod_5155(clk,rst,matrix_A[5155],matrix_B[155],mul_res1[5155]);
multi_7x28 multi_7x28_mod_5156(clk,rst,matrix_A[5156],matrix_B[156],mul_res1[5156]);
multi_7x28 multi_7x28_mod_5157(clk,rst,matrix_A[5157],matrix_B[157],mul_res1[5157]);
multi_7x28 multi_7x28_mod_5158(clk,rst,matrix_A[5158],matrix_B[158],mul_res1[5158]);
multi_7x28 multi_7x28_mod_5159(clk,rst,matrix_A[5159],matrix_B[159],mul_res1[5159]);
multi_7x28 multi_7x28_mod_5160(clk,rst,matrix_A[5160],matrix_B[160],mul_res1[5160]);
multi_7x28 multi_7x28_mod_5161(clk,rst,matrix_A[5161],matrix_B[161],mul_res1[5161]);
multi_7x28 multi_7x28_mod_5162(clk,rst,matrix_A[5162],matrix_B[162],mul_res1[5162]);
multi_7x28 multi_7x28_mod_5163(clk,rst,matrix_A[5163],matrix_B[163],mul_res1[5163]);
multi_7x28 multi_7x28_mod_5164(clk,rst,matrix_A[5164],matrix_B[164],mul_res1[5164]);
multi_7x28 multi_7x28_mod_5165(clk,rst,matrix_A[5165],matrix_B[165],mul_res1[5165]);
multi_7x28 multi_7x28_mod_5166(clk,rst,matrix_A[5166],matrix_B[166],mul_res1[5166]);
multi_7x28 multi_7x28_mod_5167(clk,rst,matrix_A[5167],matrix_B[167],mul_res1[5167]);
multi_7x28 multi_7x28_mod_5168(clk,rst,matrix_A[5168],matrix_B[168],mul_res1[5168]);
multi_7x28 multi_7x28_mod_5169(clk,rst,matrix_A[5169],matrix_B[169],mul_res1[5169]);
multi_7x28 multi_7x28_mod_5170(clk,rst,matrix_A[5170],matrix_B[170],mul_res1[5170]);
multi_7x28 multi_7x28_mod_5171(clk,rst,matrix_A[5171],matrix_B[171],mul_res1[5171]);
multi_7x28 multi_7x28_mod_5172(clk,rst,matrix_A[5172],matrix_B[172],mul_res1[5172]);
multi_7x28 multi_7x28_mod_5173(clk,rst,matrix_A[5173],matrix_B[173],mul_res1[5173]);
multi_7x28 multi_7x28_mod_5174(clk,rst,matrix_A[5174],matrix_B[174],mul_res1[5174]);
multi_7x28 multi_7x28_mod_5175(clk,rst,matrix_A[5175],matrix_B[175],mul_res1[5175]);
multi_7x28 multi_7x28_mod_5176(clk,rst,matrix_A[5176],matrix_B[176],mul_res1[5176]);
multi_7x28 multi_7x28_mod_5177(clk,rst,matrix_A[5177],matrix_B[177],mul_res1[5177]);
multi_7x28 multi_7x28_mod_5178(clk,rst,matrix_A[5178],matrix_B[178],mul_res1[5178]);
multi_7x28 multi_7x28_mod_5179(clk,rst,matrix_A[5179],matrix_B[179],mul_res1[5179]);
multi_7x28 multi_7x28_mod_5180(clk,rst,matrix_A[5180],matrix_B[180],mul_res1[5180]);
multi_7x28 multi_7x28_mod_5181(clk,rst,matrix_A[5181],matrix_B[181],mul_res1[5181]);
multi_7x28 multi_7x28_mod_5182(clk,rst,matrix_A[5182],matrix_B[182],mul_res1[5182]);
multi_7x28 multi_7x28_mod_5183(clk,rst,matrix_A[5183],matrix_B[183],mul_res1[5183]);
multi_7x28 multi_7x28_mod_5184(clk,rst,matrix_A[5184],matrix_B[184],mul_res1[5184]);
multi_7x28 multi_7x28_mod_5185(clk,rst,matrix_A[5185],matrix_B[185],mul_res1[5185]);
multi_7x28 multi_7x28_mod_5186(clk,rst,matrix_A[5186],matrix_B[186],mul_res1[5186]);
multi_7x28 multi_7x28_mod_5187(clk,rst,matrix_A[5187],matrix_B[187],mul_res1[5187]);
multi_7x28 multi_7x28_mod_5188(clk,rst,matrix_A[5188],matrix_B[188],mul_res1[5188]);
multi_7x28 multi_7x28_mod_5189(clk,rst,matrix_A[5189],matrix_B[189],mul_res1[5189]);
multi_7x28 multi_7x28_mod_5190(clk,rst,matrix_A[5190],matrix_B[190],mul_res1[5190]);
multi_7x28 multi_7x28_mod_5191(clk,rst,matrix_A[5191],matrix_B[191],mul_res1[5191]);
multi_7x28 multi_7x28_mod_5192(clk,rst,matrix_A[5192],matrix_B[192],mul_res1[5192]);
multi_7x28 multi_7x28_mod_5193(clk,rst,matrix_A[5193],matrix_B[193],mul_res1[5193]);
multi_7x28 multi_7x28_mod_5194(clk,rst,matrix_A[5194],matrix_B[194],mul_res1[5194]);
multi_7x28 multi_7x28_mod_5195(clk,rst,matrix_A[5195],matrix_B[195],mul_res1[5195]);
multi_7x28 multi_7x28_mod_5196(clk,rst,matrix_A[5196],matrix_B[196],mul_res1[5196]);
multi_7x28 multi_7x28_mod_5197(clk,rst,matrix_A[5197],matrix_B[197],mul_res1[5197]);
multi_7x28 multi_7x28_mod_5198(clk,rst,matrix_A[5198],matrix_B[198],mul_res1[5198]);
multi_7x28 multi_7x28_mod_5199(clk,rst,matrix_A[5199],matrix_B[199],mul_res1[5199]);
multi_7x28 multi_7x28_mod_5200(clk,rst,matrix_A[5200],matrix_B[0],mul_res1[5200]);
multi_7x28 multi_7x28_mod_5201(clk,rst,matrix_A[5201],matrix_B[1],mul_res1[5201]);
multi_7x28 multi_7x28_mod_5202(clk,rst,matrix_A[5202],matrix_B[2],mul_res1[5202]);
multi_7x28 multi_7x28_mod_5203(clk,rst,matrix_A[5203],matrix_B[3],mul_res1[5203]);
multi_7x28 multi_7x28_mod_5204(clk,rst,matrix_A[5204],matrix_B[4],mul_res1[5204]);
multi_7x28 multi_7x28_mod_5205(clk,rst,matrix_A[5205],matrix_B[5],mul_res1[5205]);
multi_7x28 multi_7x28_mod_5206(clk,rst,matrix_A[5206],matrix_B[6],mul_res1[5206]);
multi_7x28 multi_7x28_mod_5207(clk,rst,matrix_A[5207],matrix_B[7],mul_res1[5207]);
multi_7x28 multi_7x28_mod_5208(clk,rst,matrix_A[5208],matrix_B[8],mul_res1[5208]);
multi_7x28 multi_7x28_mod_5209(clk,rst,matrix_A[5209],matrix_B[9],mul_res1[5209]);
multi_7x28 multi_7x28_mod_5210(clk,rst,matrix_A[5210],matrix_B[10],mul_res1[5210]);
multi_7x28 multi_7x28_mod_5211(clk,rst,matrix_A[5211],matrix_B[11],mul_res1[5211]);
multi_7x28 multi_7x28_mod_5212(clk,rst,matrix_A[5212],matrix_B[12],mul_res1[5212]);
multi_7x28 multi_7x28_mod_5213(clk,rst,matrix_A[5213],matrix_B[13],mul_res1[5213]);
multi_7x28 multi_7x28_mod_5214(clk,rst,matrix_A[5214],matrix_B[14],mul_res1[5214]);
multi_7x28 multi_7x28_mod_5215(clk,rst,matrix_A[5215],matrix_B[15],mul_res1[5215]);
multi_7x28 multi_7x28_mod_5216(clk,rst,matrix_A[5216],matrix_B[16],mul_res1[5216]);
multi_7x28 multi_7x28_mod_5217(clk,rst,matrix_A[5217],matrix_B[17],mul_res1[5217]);
multi_7x28 multi_7x28_mod_5218(clk,rst,matrix_A[5218],matrix_B[18],mul_res1[5218]);
multi_7x28 multi_7x28_mod_5219(clk,rst,matrix_A[5219],matrix_B[19],mul_res1[5219]);
multi_7x28 multi_7x28_mod_5220(clk,rst,matrix_A[5220],matrix_B[20],mul_res1[5220]);
multi_7x28 multi_7x28_mod_5221(clk,rst,matrix_A[5221],matrix_B[21],mul_res1[5221]);
multi_7x28 multi_7x28_mod_5222(clk,rst,matrix_A[5222],matrix_B[22],mul_res1[5222]);
multi_7x28 multi_7x28_mod_5223(clk,rst,matrix_A[5223],matrix_B[23],mul_res1[5223]);
multi_7x28 multi_7x28_mod_5224(clk,rst,matrix_A[5224],matrix_B[24],mul_res1[5224]);
multi_7x28 multi_7x28_mod_5225(clk,rst,matrix_A[5225],matrix_B[25],mul_res1[5225]);
multi_7x28 multi_7x28_mod_5226(clk,rst,matrix_A[5226],matrix_B[26],mul_res1[5226]);
multi_7x28 multi_7x28_mod_5227(clk,rst,matrix_A[5227],matrix_B[27],mul_res1[5227]);
multi_7x28 multi_7x28_mod_5228(clk,rst,matrix_A[5228],matrix_B[28],mul_res1[5228]);
multi_7x28 multi_7x28_mod_5229(clk,rst,matrix_A[5229],matrix_B[29],mul_res1[5229]);
multi_7x28 multi_7x28_mod_5230(clk,rst,matrix_A[5230],matrix_B[30],mul_res1[5230]);
multi_7x28 multi_7x28_mod_5231(clk,rst,matrix_A[5231],matrix_B[31],mul_res1[5231]);
multi_7x28 multi_7x28_mod_5232(clk,rst,matrix_A[5232],matrix_B[32],mul_res1[5232]);
multi_7x28 multi_7x28_mod_5233(clk,rst,matrix_A[5233],matrix_B[33],mul_res1[5233]);
multi_7x28 multi_7x28_mod_5234(clk,rst,matrix_A[5234],matrix_B[34],mul_res1[5234]);
multi_7x28 multi_7x28_mod_5235(clk,rst,matrix_A[5235],matrix_B[35],mul_res1[5235]);
multi_7x28 multi_7x28_mod_5236(clk,rst,matrix_A[5236],matrix_B[36],mul_res1[5236]);
multi_7x28 multi_7x28_mod_5237(clk,rst,matrix_A[5237],matrix_B[37],mul_res1[5237]);
multi_7x28 multi_7x28_mod_5238(clk,rst,matrix_A[5238],matrix_B[38],mul_res1[5238]);
multi_7x28 multi_7x28_mod_5239(clk,rst,matrix_A[5239],matrix_B[39],mul_res1[5239]);
multi_7x28 multi_7x28_mod_5240(clk,rst,matrix_A[5240],matrix_B[40],mul_res1[5240]);
multi_7x28 multi_7x28_mod_5241(clk,rst,matrix_A[5241],matrix_B[41],mul_res1[5241]);
multi_7x28 multi_7x28_mod_5242(clk,rst,matrix_A[5242],matrix_B[42],mul_res1[5242]);
multi_7x28 multi_7x28_mod_5243(clk,rst,matrix_A[5243],matrix_B[43],mul_res1[5243]);
multi_7x28 multi_7x28_mod_5244(clk,rst,matrix_A[5244],matrix_B[44],mul_res1[5244]);
multi_7x28 multi_7x28_mod_5245(clk,rst,matrix_A[5245],matrix_B[45],mul_res1[5245]);
multi_7x28 multi_7x28_mod_5246(clk,rst,matrix_A[5246],matrix_B[46],mul_res1[5246]);
multi_7x28 multi_7x28_mod_5247(clk,rst,matrix_A[5247],matrix_B[47],mul_res1[5247]);
multi_7x28 multi_7x28_mod_5248(clk,rst,matrix_A[5248],matrix_B[48],mul_res1[5248]);
multi_7x28 multi_7x28_mod_5249(clk,rst,matrix_A[5249],matrix_B[49],mul_res1[5249]);
multi_7x28 multi_7x28_mod_5250(clk,rst,matrix_A[5250],matrix_B[50],mul_res1[5250]);
multi_7x28 multi_7x28_mod_5251(clk,rst,matrix_A[5251],matrix_B[51],mul_res1[5251]);
multi_7x28 multi_7x28_mod_5252(clk,rst,matrix_A[5252],matrix_B[52],mul_res1[5252]);
multi_7x28 multi_7x28_mod_5253(clk,rst,matrix_A[5253],matrix_B[53],mul_res1[5253]);
multi_7x28 multi_7x28_mod_5254(clk,rst,matrix_A[5254],matrix_B[54],mul_res1[5254]);
multi_7x28 multi_7x28_mod_5255(clk,rst,matrix_A[5255],matrix_B[55],mul_res1[5255]);
multi_7x28 multi_7x28_mod_5256(clk,rst,matrix_A[5256],matrix_B[56],mul_res1[5256]);
multi_7x28 multi_7x28_mod_5257(clk,rst,matrix_A[5257],matrix_B[57],mul_res1[5257]);
multi_7x28 multi_7x28_mod_5258(clk,rst,matrix_A[5258],matrix_B[58],mul_res1[5258]);
multi_7x28 multi_7x28_mod_5259(clk,rst,matrix_A[5259],matrix_B[59],mul_res1[5259]);
multi_7x28 multi_7x28_mod_5260(clk,rst,matrix_A[5260],matrix_B[60],mul_res1[5260]);
multi_7x28 multi_7x28_mod_5261(clk,rst,matrix_A[5261],matrix_B[61],mul_res1[5261]);
multi_7x28 multi_7x28_mod_5262(clk,rst,matrix_A[5262],matrix_B[62],mul_res1[5262]);
multi_7x28 multi_7x28_mod_5263(clk,rst,matrix_A[5263],matrix_B[63],mul_res1[5263]);
multi_7x28 multi_7x28_mod_5264(clk,rst,matrix_A[5264],matrix_B[64],mul_res1[5264]);
multi_7x28 multi_7x28_mod_5265(clk,rst,matrix_A[5265],matrix_B[65],mul_res1[5265]);
multi_7x28 multi_7x28_mod_5266(clk,rst,matrix_A[5266],matrix_B[66],mul_res1[5266]);
multi_7x28 multi_7x28_mod_5267(clk,rst,matrix_A[5267],matrix_B[67],mul_res1[5267]);
multi_7x28 multi_7x28_mod_5268(clk,rst,matrix_A[5268],matrix_B[68],mul_res1[5268]);
multi_7x28 multi_7x28_mod_5269(clk,rst,matrix_A[5269],matrix_B[69],mul_res1[5269]);
multi_7x28 multi_7x28_mod_5270(clk,rst,matrix_A[5270],matrix_B[70],mul_res1[5270]);
multi_7x28 multi_7x28_mod_5271(clk,rst,matrix_A[5271],matrix_B[71],mul_res1[5271]);
multi_7x28 multi_7x28_mod_5272(clk,rst,matrix_A[5272],matrix_B[72],mul_res1[5272]);
multi_7x28 multi_7x28_mod_5273(clk,rst,matrix_A[5273],matrix_B[73],mul_res1[5273]);
multi_7x28 multi_7x28_mod_5274(clk,rst,matrix_A[5274],matrix_B[74],mul_res1[5274]);
multi_7x28 multi_7x28_mod_5275(clk,rst,matrix_A[5275],matrix_B[75],mul_res1[5275]);
multi_7x28 multi_7x28_mod_5276(clk,rst,matrix_A[5276],matrix_B[76],mul_res1[5276]);
multi_7x28 multi_7x28_mod_5277(clk,rst,matrix_A[5277],matrix_B[77],mul_res1[5277]);
multi_7x28 multi_7x28_mod_5278(clk,rst,matrix_A[5278],matrix_B[78],mul_res1[5278]);
multi_7x28 multi_7x28_mod_5279(clk,rst,matrix_A[5279],matrix_B[79],mul_res1[5279]);
multi_7x28 multi_7x28_mod_5280(clk,rst,matrix_A[5280],matrix_B[80],mul_res1[5280]);
multi_7x28 multi_7x28_mod_5281(clk,rst,matrix_A[5281],matrix_B[81],mul_res1[5281]);
multi_7x28 multi_7x28_mod_5282(clk,rst,matrix_A[5282],matrix_B[82],mul_res1[5282]);
multi_7x28 multi_7x28_mod_5283(clk,rst,matrix_A[5283],matrix_B[83],mul_res1[5283]);
multi_7x28 multi_7x28_mod_5284(clk,rst,matrix_A[5284],matrix_B[84],mul_res1[5284]);
multi_7x28 multi_7x28_mod_5285(clk,rst,matrix_A[5285],matrix_B[85],mul_res1[5285]);
multi_7x28 multi_7x28_mod_5286(clk,rst,matrix_A[5286],matrix_B[86],mul_res1[5286]);
multi_7x28 multi_7x28_mod_5287(clk,rst,matrix_A[5287],matrix_B[87],mul_res1[5287]);
multi_7x28 multi_7x28_mod_5288(clk,rst,matrix_A[5288],matrix_B[88],mul_res1[5288]);
multi_7x28 multi_7x28_mod_5289(clk,rst,matrix_A[5289],matrix_B[89],mul_res1[5289]);
multi_7x28 multi_7x28_mod_5290(clk,rst,matrix_A[5290],matrix_B[90],mul_res1[5290]);
multi_7x28 multi_7x28_mod_5291(clk,rst,matrix_A[5291],matrix_B[91],mul_res1[5291]);
multi_7x28 multi_7x28_mod_5292(clk,rst,matrix_A[5292],matrix_B[92],mul_res1[5292]);
multi_7x28 multi_7x28_mod_5293(clk,rst,matrix_A[5293],matrix_B[93],mul_res1[5293]);
multi_7x28 multi_7x28_mod_5294(clk,rst,matrix_A[5294],matrix_B[94],mul_res1[5294]);
multi_7x28 multi_7x28_mod_5295(clk,rst,matrix_A[5295],matrix_B[95],mul_res1[5295]);
multi_7x28 multi_7x28_mod_5296(clk,rst,matrix_A[5296],matrix_B[96],mul_res1[5296]);
multi_7x28 multi_7x28_mod_5297(clk,rst,matrix_A[5297],matrix_B[97],mul_res1[5297]);
multi_7x28 multi_7x28_mod_5298(clk,rst,matrix_A[5298],matrix_B[98],mul_res1[5298]);
multi_7x28 multi_7x28_mod_5299(clk,rst,matrix_A[5299],matrix_B[99],mul_res1[5299]);
multi_7x28 multi_7x28_mod_5300(clk,rst,matrix_A[5300],matrix_B[100],mul_res1[5300]);
multi_7x28 multi_7x28_mod_5301(clk,rst,matrix_A[5301],matrix_B[101],mul_res1[5301]);
multi_7x28 multi_7x28_mod_5302(clk,rst,matrix_A[5302],matrix_B[102],mul_res1[5302]);
multi_7x28 multi_7x28_mod_5303(clk,rst,matrix_A[5303],matrix_B[103],mul_res1[5303]);
multi_7x28 multi_7x28_mod_5304(clk,rst,matrix_A[5304],matrix_B[104],mul_res1[5304]);
multi_7x28 multi_7x28_mod_5305(clk,rst,matrix_A[5305],matrix_B[105],mul_res1[5305]);
multi_7x28 multi_7x28_mod_5306(clk,rst,matrix_A[5306],matrix_B[106],mul_res1[5306]);
multi_7x28 multi_7x28_mod_5307(clk,rst,matrix_A[5307],matrix_B[107],mul_res1[5307]);
multi_7x28 multi_7x28_mod_5308(clk,rst,matrix_A[5308],matrix_B[108],mul_res1[5308]);
multi_7x28 multi_7x28_mod_5309(clk,rst,matrix_A[5309],matrix_B[109],mul_res1[5309]);
multi_7x28 multi_7x28_mod_5310(clk,rst,matrix_A[5310],matrix_B[110],mul_res1[5310]);
multi_7x28 multi_7x28_mod_5311(clk,rst,matrix_A[5311],matrix_B[111],mul_res1[5311]);
multi_7x28 multi_7x28_mod_5312(clk,rst,matrix_A[5312],matrix_B[112],mul_res1[5312]);
multi_7x28 multi_7x28_mod_5313(clk,rst,matrix_A[5313],matrix_B[113],mul_res1[5313]);
multi_7x28 multi_7x28_mod_5314(clk,rst,matrix_A[5314],matrix_B[114],mul_res1[5314]);
multi_7x28 multi_7x28_mod_5315(clk,rst,matrix_A[5315],matrix_B[115],mul_res1[5315]);
multi_7x28 multi_7x28_mod_5316(clk,rst,matrix_A[5316],matrix_B[116],mul_res1[5316]);
multi_7x28 multi_7x28_mod_5317(clk,rst,matrix_A[5317],matrix_B[117],mul_res1[5317]);
multi_7x28 multi_7x28_mod_5318(clk,rst,matrix_A[5318],matrix_B[118],mul_res1[5318]);
multi_7x28 multi_7x28_mod_5319(clk,rst,matrix_A[5319],matrix_B[119],mul_res1[5319]);
multi_7x28 multi_7x28_mod_5320(clk,rst,matrix_A[5320],matrix_B[120],mul_res1[5320]);
multi_7x28 multi_7x28_mod_5321(clk,rst,matrix_A[5321],matrix_B[121],mul_res1[5321]);
multi_7x28 multi_7x28_mod_5322(clk,rst,matrix_A[5322],matrix_B[122],mul_res1[5322]);
multi_7x28 multi_7x28_mod_5323(clk,rst,matrix_A[5323],matrix_B[123],mul_res1[5323]);
multi_7x28 multi_7x28_mod_5324(clk,rst,matrix_A[5324],matrix_B[124],mul_res1[5324]);
multi_7x28 multi_7x28_mod_5325(clk,rst,matrix_A[5325],matrix_B[125],mul_res1[5325]);
multi_7x28 multi_7x28_mod_5326(clk,rst,matrix_A[5326],matrix_B[126],mul_res1[5326]);
multi_7x28 multi_7x28_mod_5327(clk,rst,matrix_A[5327],matrix_B[127],mul_res1[5327]);
multi_7x28 multi_7x28_mod_5328(clk,rst,matrix_A[5328],matrix_B[128],mul_res1[5328]);
multi_7x28 multi_7x28_mod_5329(clk,rst,matrix_A[5329],matrix_B[129],mul_res1[5329]);
multi_7x28 multi_7x28_mod_5330(clk,rst,matrix_A[5330],matrix_B[130],mul_res1[5330]);
multi_7x28 multi_7x28_mod_5331(clk,rst,matrix_A[5331],matrix_B[131],mul_res1[5331]);
multi_7x28 multi_7x28_mod_5332(clk,rst,matrix_A[5332],matrix_B[132],mul_res1[5332]);
multi_7x28 multi_7x28_mod_5333(clk,rst,matrix_A[5333],matrix_B[133],mul_res1[5333]);
multi_7x28 multi_7x28_mod_5334(clk,rst,matrix_A[5334],matrix_B[134],mul_res1[5334]);
multi_7x28 multi_7x28_mod_5335(clk,rst,matrix_A[5335],matrix_B[135],mul_res1[5335]);
multi_7x28 multi_7x28_mod_5336(clk,rst,matrix_A[5336],matrix_B[136],mul_res1[5336]);
multi_7x28 multi_7x28_mod_5337(clk,rst,matrix_A[5337],matrix_B[137],mul_res1[5337]);
multi_7x28 multi_7x28_mod_5338(clk,rst,matrix_A[5338],matrix_B[138],mul_res1[5338]);
multi_7x28 multi_7x28_mod_5339(clk,rst,matrix_A[5339],matrix_B[139],mul_res1[5339]);
multi_7x28 multi_7x28_mod_5340(clk,rst,matrix_A[5340],matrix_B[140],mul_res1[5340]);
multi_7x28 multi_7x28_mod_5341(clk,rst,matrix_A[5341],matrix_B[141],mul_res1[5341]);
multi_7x28 multi_7x28_mod_5342(clk,rst,matrix_A[5342],matrix_B[142],mul_res1[5342]);
multi_7x28 multi_7x28_mod_5343(clk,rst,matrix_A[5343],matrix_B[143],mul_res1[5343]);
multi_7x28 multi_7x28_mod_5344(clk,rst,matrix_A[5344],matrix_B[144],mul_res1[5344]);
multi_7x28 multi_7x28_mod_5345(clk,rst,matrix_A[5345],matrix_B[145],mul_res1[5345]);
multi_7x28 multi_7x28_mod_5346(clk,rst,matrix_A[5346],matrix_B[146],mul_res1[5346]);
multi_7x28 multi_7x28_mod_5347(clk,rst,matrix_A[5347],matrix_B[147],mul_res1[5347]);
multi_7x28 multi_7x28_mod_5348(clk,rst,matrix_A[5348],matrix_B[148],mul_res1[5348]);
multi_7x28 multi_7x28_mod_5349(clk,rst,matrix_A[5349],matrix_B[149],mul_res1[5349]);
multi_7x28 multi_7x28_mod_5350(clk,rst,matrix_A[5350],matrix_B[150],mul_res1[5350]);
multi_7x28 multi_7x28_mod_5351(clk,rst,matrix_A[5351],matrix_B[151],mul_res1[5351]);
multi_7x28 multi_7x28_mod_5352(clk,rst,matrix_A[5352],matrix_B[152],mul_res1[5352]);
multi_7x28 multi_7x28_mod_5353(clk,rst,matrix_A[5353],matrix_B[153],mul_res1[5353]);
multi_7x28 multi_7x28_mod_5354(clk,rst,matrix_A[5354],matrix_B[154],mul_res1[5354]);
multi_7x28 multi_7x28_mod_5355(clk,rst,matrix_A[5355],matrix_B[155],mul_res1[5355]);
multi_7x28 multi_7x28_mod_5356(clk,rst,matrix_A[5356],matrix_B[156],mul_res1[5356]);
multi_7x28 multi_7x28_mod_5357(clk,rst,matrix_A[5357],matrix_B[157],mul_res1[5357]);
multi_7x28 multi_7x28_mod_5358(clk,rst,matrix_A[5358],matrix_B[158],mul_res1[5358]);
multi_7x28 multi_7x28_mod_5359(clk,rst,matrix_A[5359],matrix_B[159],mul_res1[5359]);
multi_7x28 multi_7x28_mod_5360(clk,rst,matrix_A[5360],matrix_B[160],mul_res1[5360]);
multi_7x28 multi_7x28_mod_5361(clk,rst,matrix_A[5361],matrix_B[161],mul_res1[5361]);
multi_7x28 multi_7x28_mod_5362(clk,rst,matrix_A[5362],matrix_B[162],mul_res1[5362]);
multi_7x28 multi_7x28_mod_5363(clk,rst,matrix_A[5363],matrix_B[163],mul_res1[5363]);
multi_7x28 multi_7x28_mod_5364(clk,rst,matrix_A[5364],matrix_B[164],mul_res1[5364]);
multi_7x28 multi_7x28_mod_5365(clk,rst,matrix_A[5365],matrix_B[165],mul_res1[5365]);
multi_7x28 multi_7x28_mod_5366(clk,rst,matrix_A[5366],matrix_B[166],mul_res1[5366]);
multi_7x28 multi_7x28_mod_5367(clk,rst,matrix_A[5367],matrix_B[167],mul_res1[5367]);
multi_7x28 multi_7x28_mod_5368(clk,rst,matrix_A[5368],matrix_B[168],mul_res1[5368]);
multi_7x28 multi_7x28_mod_5369(clk,rst,matrix_A[5369],matrix_B[169],mul_res1[5369]);
multi_7x28 multi_7x28_mod_5370(clk,rst,matrix_A[5370],matrix_B[170],mul_res1[5370]);
multi_7x28 multi_7x28_mod_5371(clk,rst,matrix_A[5371],matrix_B[171],mul_res1[5371]);
multi_7x28 multi_7x28_mod_5372(clk,rst,matrix_A[5372],matrix_B[172],mul_res1[5372]);
multi_7x28 multi_7x28_mod_5373(clk,rst,matrix_A[5373],matrix_B[173],mul_res1[5373]);
multi_7x28 multi_7x28_mod_5374(clk,rst,matrix_A[5374],matrix_B[174],mul_res1[5374]);
multi_7x28 multi_7x28_mod_5375(clk,rst,matrix_A[5375],matrix_B[175],mul_res1[5375]);
multi_7x28 multi_7x28_mod_5376(clk,rst,matrix_A[5376],matrix_B[176],mul_res1[5376]);
multi_7x28 multi_7x28_mod_5377(clk,rst,matrix_A[5377],matrix_B[177],mul_res1[5377]);
multi_7x28 multi_7x28_mod_5378(clk,rst,matrix_A[5378],matrix_B[178],mul_res1[5378]);
multi_7x28 multi_7x28_mod_5379(clk,rst,matrix_A[5379],matrix_B[179],mul_res1[5379]);
multi_7x28 multi_7x28_mod_5380(clk,rst,matrix_A[5380],matrix_B[180],mul_res1[5380]);
multi_7x28 multi_7x28_mod_5381(clk,rst,matrix_A[5381],matrix_B[181],mul_res1[5381]);
multi_7x28 multi_7x28_mod_5382(clk,rst,matrix_A[5382],matrix_B[182],mul_res1[5382]);
multi_7x28 multi_7x28_mod_5383(clk,rst,matrix_A[5383],matrix_B[183],mul_res1[5383]);
multi_7x28 multi_7x28_mod_5384(clk,rst,matrix_A[5384],matrix_B[184],mul_res1[5384]);
multi_7x28 multi_7x28_mod_5385(clk,rst,matrix_A[5385],matrix_B[185],mul_res1[5385]);
multi_7x28 multi_7x28_mod_5386(clk,rst,matrix_A[5386],matrix_B[186],mul_res1[5386]);
multi_7x28 multi_7x28_mod_5387(clk,rst,matrix_A[5387],matrix_B[187],mul_res1[5387]);
multi_7x28 multi_7x28_mod_5388(clk,rst,matrix_A[5388],matrix_B[188],mul_res1[5388]);
multi_7x28 multi_7x28_mod_5389(clk,rst,matrix_A[5389],matrix_B[189],mul_res1[5389]);
multi_7x28 multi_7x28_mod_5390(clk,rst,matrix_A[5390],matrix_B[190],mul_res1[5390]);
multi_7x28 multi_7x28_mod_5391(clk,rst,matrix_A[5391],matrix_B[191],mul_res1[5391]);
multi_7x28 multi_7x28_mod_5392(clk,rst,matrix_A[5392],matrix_B[192],mul_res1[5392]);
multi_7x28 multi_7x28_mod_5393(clk,rst,matrix_A[5393],matrix_B[193],mul_res1[5393]);
multi_7x28 multi_7x28_mod_5394(clk,rst,matrix_A[5394],matrix_B[194],mul_res1[5394]);
multi_7x28 multi_7x28_mod_5395(clk,rst,matrix_A[5395],matrix_B[195],mul_res1[5395]);
multi_7x28 multi_7x28_mod_5396(clk,rst,matrix_A[5396],matrix_B[196],mul_res1[5396]);
multi_7x28 multi_7x28_mod_5397(clk,rst,matrix_A[5397],matrix_B[197],mul_res1[5397]);
multi_7x28 multi_7x28_mod_5398(clk,rst,matrix_A[5398],matrix_B[198],mul_res1[5398]);
multi_7x28 multi_7x28_mod_5399(clk,rst,matrix_A[5399],matrix_B[199],mul_res1[5399]);
multi_7x28 multi_7x28_mod_5400(clk,rst,matrix_A[5400],matrix_B[0],mul_res1[5400]);
multi_7x28 multi_7x28_mod_5401(clk,rst,matrix_A[5401],matrix_B[1],mul_res1[5401]);
multi_7x28 multi_7x28_mod_5402(clk,rst,matrix_A[5402],matrix_B[2],mul_res1[5402]);
multi_7x28 multi_7x28_mod_5403(clk,rst,matrix_A[5403],matrix_B[3],mul_res1[5403]);
multi_7x28 multi_7x28_mod_5404(clk,rst,matrix_A[5404],matrix_B[4],mul_res1[5404]);
multi_7x28 multi_7x28_mod_5405(clk,rst,matrix_A[5405],matrix_B[5],mul_res1[5405]);
multi_7x28 multi_7x28_mod_5406(clk,rst,matrix_A[5406],matrix_B[6],mul_res1[5406]);
multi_7x28 multi_7x28_mod_5407(clk,rst,matrix_A[5407],matrix_B[7],mul_res1[5407]);
multi_7x28 multi_7x28_mod_5408(clk,rst,matrix_A[5408],matrix_B[8],mul_res1[5408]);
multi_7x28 multi_7x28_mod_5409(clk,rst,matrix_A[5409],matrix_B[9],mul_res1[5409]);
multi_7x28 multi_7x28_mod_5410(clk,rst,matrix_A[5410],matrix_B[10],mul_res1[5410]);
multi_7x28 multi_7x28_mod_5411(clk,rst,matrix_A[5411],matrix_B[11],mul_res1[5411]);
multi_7x28 multi_7x28_mod_5412(clk,rst,matrix_A[5412],matrix_B[12],mul_res1[5412]);
multi_7x28 multi_7x28_mod_5413(clk,rst,matrix_A[5413],matrix_B[13],mul_res1[5413]);
multi_7x28 multi_7x28_mod_5414(clk,rst,matrix_A[5414],matrix_B[14],mul_res1[5414]);
multi_7x28 multi_7x28_mod_5415(clk,rst,matrix_A[5415],matrix_B[15],mul_res1[5415]);
multi_7x28 multi_7x28_mod_5416(clk,rst,matrix_A[5416],matrix_B[16],mul_res1[5416]);
multi_7x28 multi_7x28_mod_5417(clk,rst,matrix_A[5417],matrix_B[17],mul_res1[5417]);
multi_7x28 multi_7x28_mod_5418(clk,rst,matrix_A[5418],matrix_B[18],mul_res1[5418]);
multi_7x28 multi_7x28_mod_5419(clk,rst,matrix_A[5419],matrix_B[19],mul_res1[5419]);
multi_7x28 multi_7x28_mod_5420(clk,rst,matrix_A[5420],matrix_B[20],mul_res1[5420]);
multi_7x28 multi_7x28_mod_5421(clk,rst,matrix_A[5421],matrix_B[21],mul_res1[5421]);
multi_7x28 multi_7x28_mod_5422(clk,rst,matrix_A[5422],matrix_B[22],mul_res1[5422]);
multi_7x28 multi_7x28_mod_5423(clk,rst,matrix_A[5423],matrix_B[23],mul_res1[5423]);
multi_7x28 multi_7x28_mod_5424(clk,rst,matrix_A[5424],matrix_B[24],mul_res1[5424]);
multi_7x28 multi_7x28_mod_5425(clk,rst,matrix_A[5425],matrix_B[25],mul_res1[5425]);
multi_7x28 multi_7x28_mod_5426(clk,rst,matrix_A[5426],matrix_B[26],mul_res1[5426]);
multi_7x28 multi_7x28_mod_5427(clk,rst,matrix_A[5427],matrix_B[27],mul_res1[5427]);
multi_7x28 multi_7x28_mod_5428(clk,rst,matrix_A[5428],matrix_B[28],mul_res1[5428]);
multi_7x28 multi_7x28_mod_5429(clk,rst,matrix_A[5429],matrix_B[29],mul_res1[5429]);
multi_7x28 multi_7x28_mod_5430(clk,rst,matrix_A[5430],matrix_B[30],mul_res1[5430]);
multi_7x28 multi_7x28_mod_5431(clk,rst,matrix_A[5431],matrix_B[31],mul_res1[5431]);
multi_7x28 multi_7x28_mod_5432(clk,rst,matrix_A[5432],matrix_B[32],mul_res1[5432]);
multi_7x28 multi_7x28_mod_5433(clk,rst,matrix_A[5433],matrix_B[33],mul_res1[5433]);
multi_7x28 multi_7x28_mod_5434(clk,rst,matrix_A[5434],matrix_B[34],mul_res1[5434]);
multi_7x28 multi_7x28_mod_5435(clk,rst,matrix_A[5435],matrix_B[35],mul_res1[5435]);
multi_7x28 multi_7x28_mod_5436(clk,rst,matrix_A[5436],matrix_B[36],mul_res1[5436]);
multi_7x28 multi_7x28_mod_5437(clk,rst,matrix_A[5437],matrix_B[37],mul_res1[5437]);
multi_7x28 multi_7x28_mod_5438(clk,rst,matrix_A[5438],matrix_B[38],mul_res1[5438]);
multi_7x28 multi_7x28_mod_5439(clk,rst,matrix_A[5439],matrix_B[39],mul_res1[5439]);
multi_7x28 multi_7x28_mod_5440(clk,rst,matrix_A[5440],matrix_B[40],mul_res1[5440]);
multi_7x28 multi_7x28_mod_5441(clk,rst,matrix_A[5441],matrix_B[41],mul_res1[5441]);
multi_7x28 multi_7x28_mod_5442(clk,rst,matrix_A[5442],matrix_B[42],mul_res1[5442]);
multi_7x28 multi_7x28_mod_5443(clk,rst,matrix_A[5443],matrix_B[43],mul_res1[5443]);
multi_7x28 multi_7x28_mod_5444(clk,rst,matrix_A[5444],matrix_B[44],mul_res1[5444]);
multi_7x28 multi_7x28_mod_5445(clk,rst,matrix_A[5445],matrix_B[45],mul_res1[5445]);
multi_7x28 multi_7x28_mod_5446(clk,rst,matrix_A[5446],matrix_B[46],mul_res1[5446]);
multi_7x28 multi_7x28_mod_5447(clk,rst,matrix_A[5447],matrix_B[47],mul_res1[5447]);
multi_7x28 multi_7x28_mod_5448(clk,rst,matrix_A[5448],matrix_B[48],mul_res1[5448]);
multi_7x28 multi_7x28_mod_5449(clk,rst,matrix_A[5449],matrix_B[49],mul_res1[5449]);
multi_7x28 multi_7x28_mod_5450(clk,rst,matrix_A[5450],matrix_B[50],mul_res1[5450]);
multi_7x28 multi_7x28_mod_5451(clk,rst,matrix_A[5451],matrix_B[51],mul_res1[5451]);
multi_7x28 multi_7x28_mod_5452(clk,rst,matrix_A[5452],matrix_B[52],mul_res1[5452]);
multi_7x28 multi_7x28_mod_5453(clk,rst,matrix_A[5453],matrix_B[53],mul_res1[5453]);
multi_7x28 multi_7x28_mod_5454(clk,rst,matrix_A[5454],matrix_B[54],mul_res1[5454]);
multi_7x28 multi_7x28_mod_5455(clk,rst,matrix_A[5455],matrix_B[55],mul_res1[5455]);
multi_7x28 multi_7x28_mod_5456(clk,rst,matrix_A[5456],matrix_B[56],mul_res1[5456]);
multi_7x28 multi_7x28_mod_5457(clk,rst,matrix_A[5457],matrix_B[57],mul_res1[5457]);
multi_7x28 multi_7x28_mod_5458(clk,rst,matrix_A[5458],matrix_B[58],mul_res1[5458]);
multi_7x28 multi_7x28_mod_5459(clk,rst,matrix_A[5459],matrix_B[59],mul_res1[5459]);
multi_7x28 multi_7x28_mod_5460(clk,rst,matrix_A[5460],matrix_B[60],mul_res1[5460]);
multi_7x28 multi_7x28_mod_5461(clk,rst,matrix_A[5461],matrix_B[61],mul_res1[5461]);
multi_7x28 multi_7x28_mod_5462(clk,rst,matrix_A[5462],matrix_B[62],mul_res1[5462]);
multi_7x28 multi_7x28_mod_5463(clk,rst,matrix_A[5463],matrix_B[63],mul_res1[5463]);
multi_7x28 multi_7x28_mod_5464(clk,rst,matrix_A[5464],matrix_B[64],mul_res1[5464]);
multi_7x28 multi_7x28_mod_5465(clk,rst,matrix_A[5465],matrix_B[65],mul_res1[5465]);
multi_7x28 multi_7x28_mod_5466(clk,rst,matrix_A[5466],matrix_B[66],mul_res1[5466]);
multi_7x28 multi_7x28_mod_5467(clk,rst,matrix_A[5467],matrix_B[67],mul_res1[5467]);
multi_7x28 multi_7x28_mod_5468(clk,rst,matrix_A[5468],matrix_B[68],mul_res1[5468]);
multi_7x28 multi_7x28_mod_5469(clk,rst,matrix_A[5469],matrix_B[69],mul_res1[5469]);
multi_7x28 multi_7x28_mod_5470(clk,rst,matrix_A[5470],matrix_B[70],mul_res1[5470]);
multi_7x28 multi_7x28_mod_5471(clk,rst,matrix_A[5471],matrix_B[71],mul_res1[5471]);
multi_7x28 multi_7x28_mod_5472(clk,rst,matrix_A[5472],matrix_B[72],mul_res1[5472]);
multi_7x28 multi_7x28_mod_5473(clk,rst,matrix_A[5473],matrix_B[73],mul_res1[5473]);
multi_7x28 multi_7x28_mod_5474(clk,rst,matrix_A[5474],matrix_B[74],mul_res1[5474]);
multi_7x28 multi_7x28_mod_5475(clk,rst,matrix_A[5475],matrix_B[75],mul_res1[5475]);
multi_7x28 multi_7x28_mod_5476(clk,rst,matrix_A[5476],matrix_B[76],mul_res1[5476]);
multi_7x28 multi_7x28_mod_5477(clk,rst,matrix_A[5477],matrix_B[77],mul_res1[5477]);
multi_7x28 multi_7x28_mod_5478(clk,rst,matrix_A[5478],matrix_B[78],mul_res1[5478]);
multi_7x28 multi_7x28_mod_5479(clk,rst,matrix_A[5479],matrix_B[79],mul_res1[5479]);
multi_7x28 multi_7x28_mod_5480(clk,rst,matrix_A[5480],matrix_B[80],mul_res1[5480]);
multi_7x28 multi_7x28_mod_5481(clk,rst,matrix_A[5481],matrix_B[81],mul_res1[5481]);
multi_7x28 multi_7x28_mod_5482(clk,rst,matrix_A[5482],matrix_B[82],mul_res1[5482]);
multi_7x28 multi_7x28_mod_5483(clk,rst,matrix_A[5483],matrix_B[83],mul_res1[5483]);
multi_7x28 multi_7x28_mod_5484(clk,rst,matrix_A[5484],matrix_B[84],mul_res1[5484]);
multi_7x28 multi_7x28_mod_5485(clk,rst,matrix_A[5485],matrix_B[85],mul_res1[5485]);
multi_7x28 multi_7x28_mod_5486(clk,rst,matrix_A[5486],matrix_B[86],mul_res1[5486]);
multi_7x28 multi_7x28_mod_5487(clk,rst,matrix_A[5487],matrix_B[87],mul_res1[5487]);
multi_7x28 multi_7x28_mod_5488(clk,rst,matrix_A[5488],matrix_B[88],mul_res1[5488]);
multi_7x28 multi_7x28_mod_5489(clk,rst,matrix_A[5489],matrix_B[89],mul_res1[5489]);
multi_7x28 multi_7x28_mod_5490(clk,rst,matrix_A[5490],matrix_B[90],mul_res1[5490]);
multi_7x28 multi_7x28_mod_5491(clk,rst,matrix_A[5491],matrix_B[91],mul_res1[5491]);
multi_7x28 multi_7x28_mod_5492(clk,rst,matrix_A[5492],matrix_B[92],mul_res1[5492]);
multi_7x28 multi_7x28_mod_5493(clk,rst,matrix_A[5493],matrix_B[93],mul_res1[5493]);
multi_7x28 multi_7x28_mod_5494(clk,rst,matrix_A[5494],matrix_B[94],mul_res1[5494]);
multi_7x28 multi_7x28_mod_5495(clk,rst,matrix_A[5495],matrix_B[95],mul_res1[5495]);
multi_7x28 multi_7x28_mod_5496(clk,rst,matrix_A[5496],matrix_B[96],mul_res1[5496]);
multi_7x28 multi_7x28_mod_5497(clk,rst,matrix_A[5497],matrix_B[97],mul_res1[5497]);
multi_7x28 multi_7x28_mod_5498(clk,rst,matrix_A[5498],matrix_B[98],mul_res1[5498]);
multi_7x28 multi_7x28_mod_5499(clk,rst,matrix_A[5499],matrix_B[99],mul_res1[5499]);
multi_7x28 multi_7x28_mod_5500(clk,rst,matrix_A[5500],matrix_B[100],mul_res1[5500]);
multi_7x28 multi_7x28_mod_5501(clk,rst,matrix_A[5501],matrix_B[101],mul_res1[5501]);
multi_7x28 multi_7x28_mod_5502(clk,rst,matrix_A[5502],matrix_B[102],mul_res1[5502]);
multi_7x28 multi_7x28_mod_5503(clk,rst,matrix_A[5503],matrix_B[103],mul_res1[5503]);
multi_7x28 multi_7x28_mod_5504(clk,rst,matrix_A[5504],matrix_B[104],mul_res1[5504]);
multi_7x28 multi_7x28_mod_5505(clk,rst,matrix_A[5505],matrix_B[105],mul_res1[5505]);
multi_7x28 multi_7x28_mod_5506(clk,rst,matrix_A[5506],matrix_B[106],mul_res1[5506]);
multi_7x28 multi_7x28_mod_5507(clk,rst,matrix_A[5507],matrix_B[107],mul_res1[5507]);
multi_7x28 multi_7x28_mod_5508(clk,rst,matrix_A[5508],matrix_B[108],mul_res1[5508]);
multi_7x28 multi_7x28_mod_5509(clk,rst,matrix_A[5509],matrix_B[109],mul_res1[5509]);
multi_7x28 multi_7x28_mod_5510(clk,rst,matrix_A[5510],matrix_B[110],mul_res1[5510]);
multi_7x28 multi_7x28_mod_5511(clk,rst,matrix_A[5511],matrix_B[111],mul_res1[5511]);
multi_7x28 multi_7x28_mod_5512(clk,rst,matrix_A[5512],matrix_B[112],mul_res1[5512]);
multi_7x28 multi_7x28_mod_5513(clk,rst,matrix_A[5513],matrix_B[113],mul_res1[5513]);
multi_7x28 multi_7x28_mod_5514(clk,rst,matrix_A[5514],matrix_B[114],mul_res1[5514]);
multi_7x28 multi_7x28_mod_5515(clk,rst,matrix_A[5515],matrix_B[115],mul_res1[5515]);
multi_7x28 multi_7x28_mod_5516(clk,rst,matrix_A[5516],matrix_B[116],mul_res1[5516]);
multi_7x28 multi_7x28_mod_5517(clk,rst,matrix_A[5517],matrix_B[117],mul_res1[5517]);
multi_7x28 multi_7x28_mod_5518(clk,rst,matrix_A[5518],matrix_B[118],mul_res1[5518]);
multi_7x28 multi_7x28_mod_5519(clk,rst,matrix_A[5519],matrix_B[119],mul_res1[5519]);
multi_7x28 multi_7x28_mod_5520(clk,rst,matrix_A[5520],matrix_B[120],mul_res1[5520]);
multi_7x28 multi_7x28_mod_5521(clk,rst,matrix_A[5521],matrix_B[121],mul_res1[5521]);
multi_7x28 multi_7x28_mod_5522(clk,rst,matrix_A[5522],matrix_B[122],mul_res1[5522]);
multi_7x28 multi_7x28_mod_5523(clk,rst,matrix_A[5523],matrix_B[123],mul_res1[5523]);
multi_7x28 multi_7x28_mod_5524(clk,rst,matrix_A[5524],matrix_B[124],mul_res1[5524]);
multi_7x28 multi_7x28_mod_5525(clk,rst,matrix_A[5525],matrix_B[125],mul_res1[5525]);
multi_7x28 multi_7x28_mod_5526(clk,rst,matrix_A[5526],matrix_B[126],mul_res1[5526]);
multi_7x28 multi_7x28_mod_5527(clk,rst,matrix_A[5527],matrix_B[127],mul_res1[5527]);
multi_7x28 multi_7x28_mod_5528(clk,rst,matrix_A[5528],matrix_B[128],mul_res1[5528]);
multi_7x28 multi_7x28_mod_5529(clk,rst,matrix_A[5529],matrix_B[129],mul_res1[5529]);
multi_7x28 multi_7x28_mod_5530(clk,rst,matrix_A[5530],matrix_B[130],mul_res1[5530]);
multi_7x28 multi_7x28_mod_5531(clk,rst,matrix_A[5531],matrix_B[131],mul_res1[5531]);
multi_7x28 multi_7x28_mod_5532(clk,rst,matrix_A[5532],matrix_B[132],mul_res1[5532]);
multi_7x28 multi_7x28_mod_5533(clk,rst,matrix_A[5533],matrix_B[133],mul_res1[5533]);
multi_7x28 multi_7x28_mod_5534(clk,rst,matrix_A[5534],matrix_B[134],mul_res1[5534]);
multi_7x28 multi_7x28_mod_5535(clk,rst,matrix_A[5535],matrix_B[135],mul_res1[5535]);
multi_7x28 multi_7x28_mod_5536(clk,rst,matrix_A[5536],matrix_B[136],mul_res1[5536]);
multi_7x28 multi_7x28_mod_5537(clk,rst,matrix_A[5537],matrix_B[137],mul_res1[5537]);
multi_7x28 multi_7x28_mod_5538(clk,rst,matrix_A[5538],matrix_B[138],mul_res1[5538]);
multi_7x28 multi_7x28_mod_5539(clk,rst,matrix_A[5539],matrix_B[139],mul_res1[5539]);
multi_7x28 multi_7x28_mod_5540(clk,rst,matrix_A[5540],matrix_B[140],mul_res1[5540]);
multi_7x28 multi_7x28_mod_5541(clk,rst,matrix_A[5541],matrix_B[141],mul_res1[5541]);
multi_7x28 multi_7x28_mod_5542(clk,rst,matrix_A[5542],matrix_B[142],mul_res1[5542]);
multi_7x28 multi_7x28_mod_5543(clk,rst,matrix_A[5543],matrix_B[143],mul_res1[5543]);
multi_7x28 multi_7x28_mod_5544(clk,rst,matrix_A[5544],matrix_B[144],mul_res1[5544]);
multi_7x28 multi_7x28_mod_5545(clk,rst,matrix_A[5545],matrix_B[145],mul_res1[5545]);
multi_7x28 multi_7x28_mod_5546(clk,rst,matrix_A[5546],matrix_B[146],mul_res1[5546]);
multi_7x28 multi_7x28_mod_5547(clk,rst,matrix_A[5547],matrix_B[147],mul_res1[5547]);
multi_7x28 multi_7x28_mod_5548(clk,rst,matrix_A[5548],matrix_B[148],mul_res1[5548]);
multi_7x28 multi_7x28_mod_5549(clk,rst,matrix_A[5549],matrix_B[149],mul_res1[5549]);
multi_7x28 multi_7x28_mod_5550(clk,rst,matrix_A[5550],matrix_B[150],mul_res1[5550]);
multi_7x28 multi_7x28_mod_5551(clk,rst,matrix_A[5551],matrix_B[151],mul_res1[5551]);
multi_7x28 multi_7x28_mod_5552(clk,rst,matrix_A[5552],matrix_B[152],mul_res1[5552]);
multi_7x28 multi_7x28_mod_5553(clk,rst,matrix_A[5553],matrix_B[153],mul_res1[5553]);
multi_7x28 multi_7x28_mod_5554(clk,rst,matrix_A[5554],matrix_B[154],mul_res1[5554]);
multi_7x28 multi_7x28_mod_5555(clk,rst,matrix_A[5555],matrix_B[155],mul_res1[5555]);
multi_7x28 multi_7x28_mod_5556(clk,rst,matrix_A[5556],matrix_B[156],mul_res1[5556]);
multi_7x28 multi_7x28_mod_5557(clk,rst,matrix_A[5557],matrix_B[157],mul_res1[5557]);
multi_7x28 multi_7x28_mod_5558(clk,rst,matrix_A[5558],matrix_B[158],mul_res1[5558]);
multi_7x28 multi_7x28_mod_5559(clk,rst,matrix_A[5559],matrix_B[159],mul_res1[5559]);
multi_7x28 multi_7x28_mod_5560(clk,rst,matrix_A[5560],matrix_B[160],mul_res1[5560]);
multi_7x28 multi_7x28_mod_5561(clk,rst,matrix_A[5561],matrix_B[161],mul_res1[5561]);
multi_7x28 multi_7x28_mod_5562(clk,rst,matrix_A[5562],matrix_B[162],mul_res1[5562]);
multi_7x28 multi_7x28_mod_5563(clk,rst,matrix_A[5563],matrix_B[163],mul_res1[5563]);
multi_7x28 multi_7x28_mod_5564(clk,rst,matrix_A[5564],matrix_B[164],mul_res1[5564]);
multi_7x28 multi_7x28_mod_5565(clk,rst,matrix_A[5565],matrix_B[165],mul_res1[5565]);
multi_7x28 multi_7x28_mod_5566(clk,rst,matrix_A[5566],matrix_B[166],mul_res1[5566]);
multi_7x28 multi_7x28_mod_5567(clk,rst,matrix_A[5567],matrix_B[167],mul_res1[5567]);
multi_7x28 multi_7x28_mod_5568(clk,rst,matrix_A[5568],matrix_B[168],mul_res1[5568]);
multi_7x28 multi_7x28_mod_5569(clk,rst,matrix_A[5569],matrix_B[169],mul_res1[5569]);
multi_7x28 multi_7x28_mod_5570(clk,rst,matrix_A[5570],matrix_B[170],mul_res1[5570]);
multi_7x28 multi_7x28_mod_5571(clk,rst,matrix_A[5571],matrix_B[171],mul_res1[5571]);
multi_7x28 multi_7x28_mod_5572(clk,rst,matrix_A[5572],matrix_B[172],mul_res1[5572]);
multi_7x28 multi_7x28_mod_5573(clk,rst,matrix_A[5573],matrix_B[173],mul_res1[5573]);
multi_7x28 multi_7x28_mod_5574(clk,rst,matrix_A[5574],matrix_B[174],mul_res1[5574]);
multi_7x28 multi_7x28_mod_5575(clk,rst,matrix_A[5575],matrix_B[175],mul_res1[5575]);
multi_7x28 multi_7x28_mod_5576(clk,rst,matrix_A[5576],matrix_B[176],mul_res1[5576]);
multi_7x28 multi_7x28_mod_5577(clk,rst,matrix_A[5577],matrix_B[177],mul_res1[5577]);
multi_7x28 multi_7x28_mod_5578(clk,rst,matrix_A[5578],matrix_B[178],mul_res1[5578]);
multi_7x28 multi_7x28_mod_5579(clk,rst,matrix_A[5579],matrix_B[179],mul_res1[5579]);
multi_7x28 multi_7x28_mod_5580(clk,rst,matrix_A[5580],matrix_B[180],mul_res1[5580]);
multi_7x28 multi_7x28_mod_5581(clk,rst,matrix_A[5581],matrix_B[181],mul_res1[5581]);
multi_7x28 multi_7x28_mod_5582(clk,rst,matrix_A[5582],matrix_B[182],mul_res1[5582]);
multi_7x28 multi_7x28_mod_5583(clk,rst,matrix_A[5583],matrix_B[183],mul_res1[5583]);
multi_7x28 multi_7x28_mod_5584(clk,rst,matrix_A[5584],matrix_B[184],mul_res1[5584]);
multi_7x28 multi_7x28_mod_5585(clk,rst,matrix_A[5585],matrix_B[185],mul_res1[5585]);
multi_7x28 multi_7x28_mod_5586(clk,rst,matrix_A[5586],matrix_B[186],mul_res1[5586]);
multi_7x28 multi_7x28_mod_5587(clk,rst,matrix_A[5587],matrix_B[187],mul_res1[5587]);
multi_7x28 multi_7x28_mod_5588(clk,rst,matrix_A[5588],matrix_B[188],mul_res1[5588]);
multi_7x28 multi_7x28_mod_5589(clk,rst,matrix_A[5589],matrix_B[189],mul_res1[5589]);
multi_7x28 multi_7x28_mod_5590(clk,rst,matrix_A[5590],matrix_B[190],mul_res1[5590]);
multi_7x28 multi_7x28_mod_5591(clk,rst,matrix_A[5591],matrix_B[191],mul_res1[5591]);
multi_7x28 multi_7x28_mod_5592(clk,rst,matrix_A[5592],matrix_B[192],mul_res1[5592]);
multi_7x28 multi_7x28_mod_5593(clk,rst,matrix_A[5593],matrix_B[193],mul_res1[5593]);
multi_7x28 multi_7x28_mod_5594(clk,rst,matrix_A[5594],matrix_B[194],mul_res1[5594]);
multi_7x28 multi_7x28_mod_5595(clk,rst,matrix_A[5595],matrix_B[195],mul_res1[5595]);
multi_7x28 multi_7x28_mod_5596(clk,rst,matrix_A[5596],matrix_B[196],mul_res1[5596]);
multi_7x28 multi_7x28_mod_5597(clk,rst,matrix_A[5597],matrix_B[197],mul_res1[5597]);
multi_7x28 multi_7x28_mod_5598(clk,rst,matrix_A[5598],matrix_B[198],mul_res1[5598]);
multi_7x28 multi_7x28_mod_5599(clk,rst,matrix_A[5599],matrix_B[199],mul_res1[5599]);
multi_7x28 multi_7x28_mod_5600(clk,rst,matrix_A[5600],matrix_B[0],mul_res1[5600]);
multi_7x28 multi_7x28_mod_5601(clk,rst,matrix_A[5601],matrix_B[1],mul_res1[5601]);
multi_7x28 multi_7x28_mod_5602(clk,rst,matrix_A[5602],matrix_B[2],mul_res1[5602]);
multi_7x28 multi_7x28_mod_5603(clk,rst,matrix_A[5603],matrix_B[3],mul_res1[5603]);
multi_7x28 multi_7x28_mod_5604(clk,rst,matrix_A[5604],matrix_B[4],mul_res1[5604]);
multi_7x28 multi_7x28_mod_5605(clk,rst,matrix_A[5605],matrix_B[5],mul_res1[5605]);
multi_7x28 multi_7x28_mod_5606(clk,rst,matrix_A[5606],matrix_B[6],mul_res1[5606]);
multi_7x28 multi_7x28_mod_5607(clk,rst,matrix_A[5607],matrix_B[7],mul_res1[5607]);
multi_7x28 multi_7x28_mod_5608(clk,rst,matrix_A[5608],matrix_B[8],mul_res1[5608]);
multi_7x28 multi_7x28_mod_5609(clk,rst,matrix_A[5609],matrix_B[9],mul_res1[5609]);
multi_7x28 multi_7x28_mod_5610(clk,rst,matrix_A[5610],matrix_B[10],mul_res1[5610]);
multi_7x28 multi_7x28_mod_5611(clk,rst,matrix_A[5611],matrix_B[11],mul_res1[5611]);
multi_7x28 multi_7x28_mod_5612(clk,rst,matrix_A[5612],matrix_B[12],mul_res1[5612]);
multi_7x28 multi_7x28_mod_5613(clk,rst,matrix_A[5613],matrix_B[13],mul_res1[5613]);
multi_7x28 multi_7x28_mod_5614(clk,rst,matrix_A[5614],matrix_B[14],mul_res1[5614]);
multi_7x28 multi_7x28_mod_5615(clk,rst,matrix_A[5615],matrix_B[15],mul_res1[5615]);
multi_7x28 multi_7x28_mod_5616(clk,rst,matrix_A[5616],matrix_B[16],mul_res1[5616]);
multi_7x28 multi_7x28_mod_5617(clk,rst,matrix_A[5617],matrix_B[17],mul_res1[5617]);
multi_7x28 multi_7x28_mod_5618(clk,rst,matrix_A[5618],matrix_B[18],mul_res1[5618]);
multi_7x28 multi_7x28_mod_5619(clk,rst,matrix_A[5619],matrix_B[19],mul_res1[5619]);
multi_7x28 multi_7x28_mod_5620(clk,rst,matrix_A[5620],matrix_B[20],mul_res1[5620]);
multi_7x28 multi_7x28_mod_5621(clk,rst,matrix_A[5621],matrix_B[21],mul_res1[5621]);
multi_7x28 multi_7x28_mod_5622(clk,rst,matrix_A[5622],matrix_B[22],mul_res1[5622]);
multi_7x28 multi_7x28_mod_5623(clk,rst,matrix_A[5623],matrix_B[23],mul_res1[5623]);
multi_7x28 multi_7x28_mod_5624(clk,rst,matrix_A[5624],matrix_B[24],mul_res1[5624]);
multi_7x28 multi_7x28_mod_5625(clk,rst,matrix_A[5625],matrix_B[25],mul_res1[5625]);
multi_7x28 multi_7x28_mod_5626(clk,rst,matrix_A[5626],matrix_B[26],mul_res1[5626]);
multi_7x28 multi_7x28_mod_5627(clk,rst,matrix_A[5627],matrix_B[27],mul_res1[5627]);
multi_7x28 multi_7x28_mod_5628(clk,rst,matrix_A[5628],matrix_B[28],mul_res1[5628]);
multi_7x28 multi_7x28_mod_5629(clk,rst,matrix_A[5629],matrix_B[29],mul_res1[5629]);
multi_7x28 multi_7x28_mod_5630(clk,rst,matrix_A[5630],matrix_B[30],mul_res1[5630]);
multi_7x28 multi_7x28_mod_5631(clk,rst,matrix_A[5631],matrix_B[31],mul_res1[5631]);
multi_7x28 multi_7x28_mod_5632(clk,rst,matrix_A[5632],matrix_B[32],mul_res1[5632]);
multi_7x28 multi_7x28_mod_5633(clk,rst,matrix_A[5633],matrix_B[33],mul_res1[5633]);
multi_7x28 multi_7x28_mod_5634(clk,rst,matrix_A[5634],matrix_B[34],mul_res1[5634]);
multi_7x28 multi_7x28_mod_5635(clk,rst,matrix_A[5635],matrix_B[35],mul_res1[5635]);
multi_7x28 multi_7x28_mod_5636(clk,rst,matrix_A[5636],matrix_B[36],mul_res1[5636]);
multi_7x28 multi_7x28_mod_5637(clk,rst,matrix_A[5637],matrix_B[37],mul_res1[5637]);
multi_7x28 multi_7x28_mod_5638(clk,rst,matrix_A[5638],matrix_B[38],mul_res1[5638]);
multi_7x28 multi_7x28_mod_5639(clk,rst,matrix_A[5639],matrix_B[39],mul_res1[5639]);
multi_7x28 multi_7x28_mod_5640(clk,rst,matrix_A[5640],matrix_B[40],mul_res1[5640]);
multi_7x28 multi_7x28_mod_5641(clk,rst,matrix_A[5641],matrix_B[41],mul_res1[5641]);
multi_7x28 multi_7x28_mod_5642(clk,rst,matrix_A[5642],matrix_B[42],mul_res1[5642]);
multi_7x28 multi_7x28_mod_5643(clk,rst,matrix_A[5643],matrix_B[43],mul_res1[5643]);
multi_7x28 multi_7x28_mod_5644(clk,rst,matrix_A[5644],matrix_B[44],mul_res1[5644]);
multi_7x28 multi_7x28_mod_5645(clk,rst,matrix_A[5645],matrix_B[45],mul_res1[5645]);
multi_7x28 multi_7x28_mod_5646(clk,rst,matrix_A[5646],matrix_B[46],mul_res1[5646]);
multi_7x28 multi_7x28_mod_5647(clk,rst,matrix_A[5647],matrix_B[47],mul_res1[5647]);
multi_7x28 multi_7x28_mod_5648(clk,rst,matrix_A[5648],matrix_B[48],mul_res1[5648]);
multi_7x28 multi_7x28_mod_5649(clk,rst,matrix_A[5649],matrix_B[49],mul_res1[5649]);
multi_7x28 multi_7x28_mod_5650(clk,rst,matrix_A[5650],matrix_B[50],mul_res1[5650]);
multi_7x28 multi_7x28_mod_5651(clk,rst,matrix_A[5651],matrix_B[51],mul_res1[5651]);
multi_7x28 multi_7x28_mod_5652(clk,rst,matrix_A[5652],matrix_B[52],mul_res1[5652]);
multi_7x28 multi_7x28_mod_5653(clk,rst,matrix_A[5653],matrix_B[53],mul_res1[5653]);
multi_7x28 multi_7x28_mod_5654(clk,rst,matrix_A[5654],matrix_B[54],mul_res1[5654]);
multi_7x28 multi_7x28_mod_5655(clk,rst,matrix_A[5655],matrix_B[55],mul_res1[5655]);
multi_7x28 multi_7x28_mod_5656(clk,rst,matrix_A[5656],matrix_B[56],mul_res1[5656]);
multi_7x28 multi_7x28_mod_5657(clk,rst,matrix_A[5657],matrix_B[57],mul_res1[5657]);
multi_7x28 multi_7x28_mod_5658(clk,rst,matrix_A[5658],matrix_B[58],mul_res1[5658]);
multi_7x28 multi_7x28_mod_5659(clk,rst,matrix_A[5659],matrix_B[59],mul_res1[5659]);
multi_7x28 multi_7x28_mod_5660(clk,rst,matrix_A[5660],matrix_B[60],mul_res1[5660]);
multi_7x28 multi_7x28_mod_5661(clk,rst,matrix_A[5661],matrix_B[61],mul_res1[5661]);
multi_7x28 multi_7x28_mod_5662(clk,rst,matrix_A[5662],matrix_B[62],mul_res1[5662]);
multi_7x28 multi_7x28_mod_5663(clk,rst,matrix_A[5663],matrix_B[63],mul_res1[5663]);
multi_7x28 multi_7x28_mod_5664(clk,rst,matrix_A[5664],matrix_B[64],mul_res1[5664]);
multi_7x28 multi_7x28_mod_5665(clk,rst,matrix_A[5665],matrix_B[65],mul_res1[5665]);
multi_7x28 multi_7x28_mod_5666(clk,rst,matrix_A[5666],matrix_B[66],mul_res1[5666]);
multi_7x28 multi_7x28_mod_5667(clk,rst,matrix_A[5667],matrix_B[67],mul_res1[5667]);
multi_7x28 multi_7x28_mod_5668(clk,rst,matrix_A[5668],matrix_B[68],mul_res1[5668]);
multi_7x28 multi_7x28_mod_5669(clk,rst,matrix_A[5669],matrix_B[69],mul_res1[5669]);
multi_7x28 multi_7x28_mod_5670(clk,rst,matrix_A[5670],matrix_B[70],mul_res1[5670]);
multi_7x28 multi_7x28_mod_5671(clk,rst,matrix_A[5671],matrix_B[71],mul_res1[5671]);
multi_7x28 multi_7x28_mod_5672(clk,rst,matrix_A[5672],matrix_B[72],mul_res1[5672]);
multi_7x28 multi_7x28_mod_5673(clk,rst,matrix_A[5673],matrix_B[73],mul_res1[5673]);
multi_7x28 multi_7x28_mod_5674(clk,rst,matrix_A[5674],matrix_B[74],mul_res1[5674]);
multi_7x28 multi_7x28_mod_5675(clk,rst,matrix_A[5675],matrix_B[75],mul_res1[5675]);
multi_7x28 multi_7x28_mod_5676(clk,rst,matrix_A[5676],matrix_B[76],mul_res1[5676]);
multi_7x28 multi_7x28_mod_5677(clk,rst,matrix_A[5677],matrix_B[77],mul_res1[5677]);
multi_7x28 multi_7x28_mod_5678(clk,rst,matrix_A[5678],matrix_B[78],mul_res1[5678]);
multi_7x28 multi_7x28_mod_5679(clk,rst,matrix_A[5679],matrix_B[79],mul_res1[5679]);
multi_7x28 multi_7x28_mod_5680(clk,rst,matrix_A[5680],matrix_B[80],mul_res1[5680]);
multi_7x28 multi_7x28_mod_5681(clk,rst,matrix_A[5681],matrix_B[81],mul_res1[5681]);
multi_7x28 multi_7x28_mod_5682(clk,rst,matrix_A[5682],matrix_B[82],mul_res1[5682]);
multi_7x28 multi_7x28_mod_5683(clk,rst,matrix_A[5683],matrix_B[83],mul_res1[5683]);
multi_7x28 multi_7x28_mod_5684(clk,rst,matrix_A[5684],matrix_B[84],mul_res1[5684]);
multi_7x28 multi_7x28_mod_5685(clk,rst,matrix_A[5685],matrix_B[85],mul_res1[5685]);
multi_7x28 multi_7x28_mod_5686(clk,rst,matrix_A[5686],matrix_B[86],mul_res1[5686]);
multi_7x28 multi_7x28_mod_5687(clk,rst,matrix_A[5687],matrix_B[87],mul_res1[5687]);
multi_7x28 multi_7x28_mod_5688(clk,rst,matrix_A[5688],matrix_B[88],mul_res1[5688]);
multi_7x28 multi_7x28_mod_5689(clk,rst,matrix_A[5689],matrix_B[89],mul_res1[5689]);
multi_7x28 multi_7x28_mod_5690(clk,rst,matrix_A[5690],matrix_B[90],mul_res1[5690]);
multi_7x28 multi_7x28_mod_5691(clk,rst,matrix_A[5691],matrix_B[91],mul_res1[5691]);
multi_7x28 multi_7x28_mod_5692(clk,rst,matrix_A[5692],matrix_B[92],mul_res1[5692]);
multi_7x28 multi_7x28_mod_5693(clk,rst,matrix_A[5693],matrix_B[93],mul_res1[5693]);
multi_7x28 multi_7x28_mod_5694(clk,rst,matrix_A[5694],matrix_B[94],mul_res1[5694]);
multi_7x28 multi_7x28_mod_5695(clk,rst,matrix_A[5695],matrix_B[95],mul_res1[5695]);
multi_7x28 multi_7x28_mod_5696(clk,rst,matrix_A[5696],matrix_B[96],mul_res1[5696]);
multi_7x28 multi_7x28_mod_5697(clk,rst,matrix_A[5697],matrix_B[97],mul_res1[5697]);
multi_7x28 multi_7x28_mod_5698(clk,rst,matrix_A[5698],matrix_B[98],mul_res1[5698]);
multi_7x28 multi_7x28_mod_5699(clk,rst,matrix_A[5699],matrix_B[99],mul_res1[5699]);
multi_7x28 multi_7x28_mod_5700(clk,rst,matrix_A[5700],matrix_B[100],mul_res1[5700]);
multi_7x28 multi_7x28_mod_5701(clk,rst,matrix_A[5701],matrix_B[101],mul_res1[5701]);
multi_7x28 multi_7x28_mod_5702(clk,rst,matrix_A[5702],matrix_B[102],mul_res1[5702]);
multi_7x28 multi_7x28_mod_5703(clk,rst,matrix_A[5703],matrix_B[103],mul_res1[5703]);
multi_7x28 multi_7x28_mod_5704(clk,rst,matrix_A[5704],matrix_B[104],mul_res1[5704]);
multi_7x28 multi_7x28_mod_5705(clk,rst,matrix_A[5705],matrix_B[105],mul_res1[5705]);
multi_7x28 multi_7x28_mod_5706(clk,rst,matrix_A[5706],matrix_B[106],mul_res1[5706]);
multi_7x28 multi_7x28_mod_5707(clk,rst,matrix_A[5707],matrix_B[107],mul_res1[5707]);
multi_7x28 multi_7x28_mod_5708(clk,rst,matrix_A[5708],matrix_B[108],mul_res1[5708]);
multi_7x28 multi_7x28_mod_5709(clk,rst,matrix_A[5709],matrix_B[109],mul_res1[5709]);
multi_7x28 multi_7x28_mod_5710(clk,rst,matrix_A[5710],matrix_B[110],mul_res1[5710]);
multi_7x28 multi_7x28_mod_5711(clk,rst,matrix_A[5711],matrix_B[111],mul_res1[5711]);
multi_7x28 multi_7x28_mod_5712(clk,rst,matrix_A[5712],matrix_B[112],mul_res1[5712]);
multi_7x28 multi_7x28_mod_5713(clk,rst,matrix_A[5713],matrix_B[113],mul_res1[5713]);
multi_7x28 multi_7x28_mod_5714(clk,rst,matrix_A[5714],matrix_B[114],mul_res1[5714]);
multi_7x28 multi_7x28_mod_5715(clk,rst,matrix_A[5715],matrix_B[115],mul_res1[5715]);
multi_7x28 multi_7x28_mod_5716(clk,rst,matrix_A[5716],matrix_B[116],mul_res1[5716]);
multi_7x28 multi_7x28_mod_5717(clk,rst,matrix_A[5717],matrix_B[117],mul_res1[5717]);
multi_7x28 multi_7x28_mod_5718(clk,rst,matrix_A[5718],matrix_B[118],mul_res1[5718]);
multi_7x28 multi_7x28_mod_5719(clk,rst,matrix_A[5719],matrix_B[119],mul_res1[5719]);
multi_7x28 multi_7x28_mod_5720(clk,rst,matrix_A[5720],matrix_B[120],mul_res1[5720]);
multi_7x28 multi_7x28_mod_5721(clk,rst,matrix_A[5721],matrix_B[121],mul_res1[5721]);
multi_7x28 multi_7x28_mod_5722(clk,rst,matrix_A[5722],matrix_B[122],mul_res1[5722]);
multi_7x28 multi_7x28_mod_5723(clk,rst,matrix_A[5723],matrix_B[123],mul_res1[5723]);
multi_7x28 multi_7x28_mod_5724(clk,rst,matrix_A[5724],matrix_B[124],mul_res1[5724]);
multi_7x28 multi_7x28_mod_5725(clk,rst,matrix_A[5725],matrix_B[125],mul_res1[5725]);
multi_7x28 multi_7x28_mod_5726(clk,rst,matrix_A[5726],matrix_B[126],mul_res1[5726]);
multi_7x28 multi_7x28_mod_5727(clk,rst,matrix_A[5727],matrix_B[127],mul_res1[5727]);
multi_7x28 multi_7x28_mod_5728(clk,rst,matrix_A[5728],matrix_B[128],mul_res1[5728]);
multi_7x28 multi_7x28_mod_5729(clk,rst,matrix_A[5729],matrix_B[129],mul_res1[5729]);
multi_7x28 multi_7x28_mod_5730(clk,rst,matrix_A[5730],matrix_B[130],mul_res1[5730]);
multi_7x28 multi_7x28_mod_5731(clk,rst,matrix_A[5731],matrix_B[131],mul_res1[5731]);
multi_7x28 multi_7x28_mod_5732(clk,rst,matrix_A[5732],matrix_B[132],mul_res1[5732]);
multi_7x28 multi_7x28_mod_5733(clk,rst,matrix_A[5733],matrix_B[133],mul_res1[5733]);
multi_7x28 multi_7x28_mod_5734(clk,rst,matrix_A[5734],matrix_B[134],mul_res1[5734]);
multi_7x28 multi_7x28_mod_5735(clk,rst,matrix_A[5735],matrix_B[135],mul_res1[5735]);
multi_7x28 multi_7x28_mod_5736(clk,rst,matrix_A[5736],matrix_B[136],mul_res1[5736]);
multi_7x28 multi_7x28_mod_5737(clk,rst,matrix_A[5737],matrix_B[137],mul_res1[5737]);
multi_7x28 multi_7x28_mod_5738(clk,rst,matrix_A[5738],matrix_B[138],mul_res1[5738]);
multi_7x28 multi_7x28_mod_5739(clk,rst,matrix_A[5739],matrix_B[139],mul_res1[5739]);
multi_7x28 multi_7x28_mod_5740(clk,rst,matrix_A[5740],matrix_B[140],mul_res1[5740]);
multi_7x28 multi_7x28_mod_5741(clk,rst,matrix_A[5741],matrix_B[141],mul_res1[5741]);
multi_7x28 multi_7x28_mod_5742(clk,rst,matrix_A[5742],matrix_B[142],mul_res1[5742]);
multi_7x28 multi_7x28_mod_5743(clk,rst,matrix_A[5743],matrix_B[143],mul_res1[5743]);
multi_7x28 multi_7x28_mod_5744(clk,rst,matrix_A[5744],matrix_B[144],mul_res1[5744]);
multi_7x28 multi_7x28_mod_5745(clk,rst,matrix_A[5745],matrix_B[145],mul_res1[5745]);
multi_7x28 multi_7x28_mod_5746(clk,rst,matrix_A[5746],matrix_B[146],mul_res1[5746]);
multi_7x28 multi_7x28_mod_5747(clk,rst,matrix_A[5747],matrix_B[147],mul_res1[5747]);
multi_7x28 multi_7x28_mod_5748(clk,rst,matrix_A[5748],matrix_B[148],mul_res1[5748]);
multi_7x28 multi_7x28_mod_5749(clk,rst,matrix_A[5749],matrix_B[149],mul_res1[5749]);
multi_7x28 multi_7x28_mod_5750(clk,rst,matrix_A[5750],matrix_B[150],mul_res1[5750]);
multi_7x28 multi_7x28_mod_5751(clk,rst,matrix_A[5751],matrix_B[151],mul_res1[5751]);
multi_7x28 multi_7x28_mod_5752(clk,rst,matrix_A[5752],matrix_B[152],mul_res1[5752]);
multi_7x28 multi_7x28_mod_5753(clk,rst,matrix_A[5753],matrix_B[153],mul_res1[5753]);
multi_7x28 multi_7x28_mod_5754(clk,rst,matrix_A[5754],matrix_B[154],mul_res1[5754]);
multi_7x28 multi_7x28_mod_5755(clk,rst,matrix_A[5755],matrix_B[155],mul_res1[5755]);
multi_7x28 multi_7x28_mod_5756(clk,rst,matrix_A[5756],matrix_B[156],mul_res1[5756]);
multi_7x28 multi_7x28_mod_5757(clk,rst,matrix_A[5757],matrix_B[157],mul_res1[5757]);
multi_7x28 multi_7x28_mod_5758(clk,rst,matrix_A[5758],matrix_B[158],mul_res1[5758]);
multi_7x28 multi_7x28_mod_5759(clk,rst,matrix_A[5759],matrix_B[159],mul_res1[5759]);
multi_7x28 multi_7x28_mod_5760(clk,rst,matrix_A[5760],matrix_B[160],mul_res1[5760]);
multi_7x28 multi_7x28_mod_5761(clk,rst,matrix_A[5761],matrix_B[161],mul_res1[5761]);
multi_7x28 multi_7x28_mod_5762(clk,rst,matrix_A[5762],matrix_B[162],mul_res1[5762]);
multi_7x28 multi_7x28_mod_5763(clk,rst,matrix_A[5763],matrix_B[163],mul_res1[5763]);
multi_7x28 multi_7x28_mod_5764(clk,rst,matrix_A[5764],matrix_B[164],mul_res1[5764]);
multi_7x28 multi_7x28_mod_5765(clk,rst,matrix_A[5765],matrix_B[165],mul_res1[5765]);
multi_7x28 multi_7x28_mod_5766(clk,rst,matrix_A[5766],matrix_B[166],mul_res1[5766]);
multi_7x28 multi_7x28_mod_5767(clk,rst,matrix_A[5767],matrix_B[167],mul_res1[5767]);
multi_7x28 multi_7x28_mod_5768(clk,rst,matrix_A[5768],matrix_B[168],mul_res1[5768]);
multi_7x28 multi_7x28_mod_5769(clk,rst,matrix_A[5769],matrix_B[169],mul_res1[5769]);
multi_7x28 multi_7x28_mod_5770(clk,rst,matrix_A[5770],matrix_B[170],mul_res1[5770]);
multi_7x28 multi_7x28_mod_5771(clk,rst,matrix_A[5771],matrix_B[171],mul_res1[5771]);
multi_7x28 multi_7x28_mod_5772(clk,rst,matrix_A[5772],matrix_B[172],mul_res1[5772]);
multi_7x28 multi_7x28_mod_5773(clk,rst,matrix_A[5773],matrix_B[173],mul_res1[5773]);
multi_7x28 multi_7x28_mod_5774(clk,rst,matrix_A[5774],matrix_B[174],mul_res1[5774]);
multi_7x28 multi_7x28_mod_5775(clk,rst,matrix_A[5775],matrix_B[175],mul_res1[5775]);
multi_7x28 multi_7x28_mod_5776(clk,rst,matrix_A[5776],matrix_B[176],mul_res1[5776]);
multi_7x28 multi_7x28_mod_5777(clk,rst,matrix_A[5777],matrix_B[177],mul_res1[5777]);
multi_7x28 multi_7x28_mod_5778(clk,rst,matrix_A[5778],matrix_B[178],mul_res1[5778]);
multi_7x28 multi_7x28_mod_5779(clk,rst,matrix_A[5779],matrix_B[179],mul_res1[5779]);
multi_7x28 multi_7x28_mod_5780(clk,rst,matrix_A[5780],matrix_B[180],mul_res1[5780]);
multi_7x28 multi_7x28_mod_5781(clk,rst,matrix_A[5781],matrix_B[181],mul_res1[5781]);
multi_7x28 multi_7x28_mod_5782(clk,rst,matrix_A[5782],matrix_B[182],mul_res1[5782]);
multi_7x28 multi_7x28_mod_5783(clk,rst,matrix_A[5783],matrix_B[183],mul_res1[5783]);
multi_7x28 multi_7x28_mod_5784(clk,rst,matrix_A[5784],matrix_B[184],mul_res1[5784]);
multi_7x28 multi_7x28_mod_5785(clk,rst,matrix_A[5785],matrix_B[185],mul_res1[5785]);
multi_7x28 multi_7x28_mod_5786(clk,rst,matrix_A[5786],matrix_B[186],mul_res1[5786]);
multi_7x28 multi_7x28_mod_5787(clk,rst,matrix_A[5787],matrix_B[187],mul_res1[5787]);
multi_7x28 multi_7x28_mod_5788(clk,rst,matrix_A[5788],matrix_B[188],mul_res1[5788]);
multi_7x28 multi_7x28_mod_5789(clk,rst,matrix_A[5789],matrix_B[189],mul_res1[5789]);
multi_7x28 multi_7x28_mod_5790(clk,rst,matrix_A[5790],matrix_B[190],mul_res1[5790]);
multi_7x28 multi_7x28_mod_5791(clk,rst,matrix_A[5791],matrix_B[191],mul_res1[5791]);
multi_7x28 multi_7x28_mod_5792(clk,rst,matrix_A[5792],matrix_B[192],mul_res1[5792]);
multi_7x28 multi_7x28_mod_5793(clk,rst,matrix_A[5793],matrix_B[193],mul_res1[5793]);
multi_7x28 multi_7x28_mod_5794(clk,rst,matrix_A[5794],matrix_B[194],mul_res1[5794]);
multi_7x28 multi_7x28_mod_5795(clk,rst,matrix_A[5795],matrix_B[195],mul_res1[5795]);
multi_7x28 multi_7x28_mod_5796(clk,rst,matrix_A[5796],matrix_B[196],mul_res1[5796]);
multi_7x28 multi_7x28_mod_5797(clk,rst,matrix_A[5797],matrix_B[197],mul_res1[5797]);
multi_7x28 multi_7x28_mod_5798(clk,rst,matrix_A[5798],matrix_B[198],mul_res1[5798]);
multi_7x28 multi_7x28_mod_5799(clk,rst,matrix_A[5799],matrix_B[199],mul_res1[5799]);
multi_7x28 multi_7x28_mod_5800(clk,rst,matrix_A[5800],matrix_B[0],mul_res1[5800]);
multi_7x28 multi_7x28_mod_5801(clk,rst,matrix_A[5801],matrix_B[1],mul_res1[5801]);
multi_7x28 multi_7x28_mod_5802(clk,rst,matrix_A[5802],matrix_B[2],mul_res1[5802]);
multi_7x28 multi_7x28_mod_5803(clk,rst,matrix_A[5803],matrix_B[3],mul_res1[5803]);
multi_7x28 multi_7x28_mod_5804(clk,rst,matrix_A[5804],matrix_B[4],mul_res1[5804]);
multi_7x28 multi_7x28_mod_5805(clk,rst,matrix_A[5805],matrix_B[5],mul_res1[5805]);
multi_7x28 multi_7x28_mod_5806(clk,rst,matrix_A[5806],matrix_B[6],mul_res1[5806]);
multi_7x28 multi_7x28_mod_5807(clk,rst,matrix_A[5807],matrix_B[7],mul_res1[5807]);
multi_7x28 multi_7x28_mod_5808(clk,rst,matrix_A[5808],matrix_B[8],mul_res1[5808]);
multi_7x28 multi_7x28_mod_5809(clk,rst,matrix_A[5809],matrix_B[9],mul_res1[5809]);
multi_7x28 multi_7x28_mod_5810(clk,rst,matrix_A[5810],matrix_B[10],mul_res1[5810]);
multi_7x28 multi_7x28_mod_5811(clk,rst,matrix_A[5811],matrix_B[11],mul_res1[5811]);
multi_7x28 multi_7x28_mod_5812(clk,rst,matrix_A[5812],matrix_B[12],mul_res1[5812]);
multi_7x28 multi_7x28_mod_5813(clk,rst,matrix_A[5813],matrix_B[13],mul_res1[5813]);
multi_7x28 multi_7x28_mod_5814(clk,rst,matrix_A[5814],matrix_B[14],mul_res1[5814]);
multi_7x28 multi_7x28_mod_5815(clk,rst,matrix_A[5815],matrix_B[15],mul_res1[5815]);
multi_7x28 multi_7x28_mod_5816(clk,rst,matrix_A[5816],matrix_B[16],mul_res1[5816]);
multi_7x28 multi_7x28_mod_5817(clk,rst,matrix_A[5817],matrix_B[17],mul_res1[5817]);
multi_7x28 multi_7x28_mod_5818(clk,rst,matrix_A[5818],matrix_B[18],mul_res1[5818]);
multi_7x28 multi_7x28_mod_5819(clk,rst,matrix_A[5819],matrix_B[19],mul_res1[5819]);
multi_7x28 multi_7x28_mod_5820(clk,rst,matrix_A[5820],matrix_B[20],mul_res1[5820]);
multi_7x28 multi_7x28_mod_5821(clk,rst,matrix_A[5821],matrix_B[21],mul_res1[5821]);
multi_7x28 multi_7x28_mod_5822(clk,rst,matrix_A[5822],matrix_B[22],mul_res1[5822]);
multi_7x28 multi_7x28_mod_5823(clk,rst,matrix_A[5823],matrix_B[23],mul_res1[5823]);
multi_7x28 multi_7x28_mod_5824(clk,rst,matrix_A[5824],matrix_B[24],mul_res1[5824]);
multi_7x28 multi_7x28_mod_5825(clk,rst,matrix_A[5825],matrix_B[25],mul_res1[5825]);
multi_7x28 multi_7x28_mod_5826(clk,rst,matrix_A[5826],matrix_B[26],mul_res1[5826]);
multi_7x28 multi_7x28_mod_5827(clk,rst,matrix_A[5827],matrix_B[27],mul_res1[5827]);
multi_7x28 multi_7x28_mod_5828(clk,rst,matrix_A[5828],matrix_B[28],mul_res1[5828]);
multi_7x28 multi_7x28_mod_5829(clk,rst,matrix_A[5829],matrix_B[29],mul_res1[5829]);
multi_7x28 multi_7x28_mod_5830(clk,rst,matrix_A[5830],matrix_B[30],mul_res1[5830]);
multi_7x28 multi_7x28_mod_5831(clk,rst,matrix_A[5831],matrix_B[31],mul_res1[5831]);
multi_7x28 multi_7x28_mod_5832(clk,rst,matrix_A[5832],matrix_B[32],mul_res1[5832]);
multi_7x28 multi_7x28_mod_5833(clk,rst,matrix_A[5833],matrix_B[33],mul_res1[5833]);
multi_7x28 multi_7x28_mod_5834(clk,rst,matrix_A[5834],matrix_B[34],mul_res1[5834]);
multi_7x28 multi_7x28_mod_5835(clk,rst,matrix_A[5835],matrix_B[35],mul_res1[5835]);
multi_7x28 multi_7x28_mod_5836(clk,rst,matrix_A[5836],matrix_B[36],mul_res1[5836]);
multi_7x28 multi_7x28_mod_5837(clk,rst,matrix_A[5837],matrix_B[37],mul_res1[5837]);
multi_7x28 multi_7x28_mod_5838(clk,rst,matrix_A[5838],matrix_B[38],mul_res1[5838]);
multi_7x28 multi_7x28_mod_5839(clk,rst,matrix_A[5839],matrix_B[39],mul_res1[5839]);
multi_7x28 multi_7x28_mod_5840(clk,rst,matrix_A[5840],matrix_B[40],mul_res1[5840]);
multi_7x28 multi_7x28_mod_5841(clk,rst,matrix_A[5841],matrix_B[41],mul_res1[5841]);
multi_7x28 multi_7x28_mod_5842(clk,rst,matrix_A[5842],matrix_B[42],mul_res1[5842]);
multi_7x28 multi_7x28_mod_5843(clk,rst,matrix_A[5843],matrix_B[43],mul_res1[5843]);
multi_7x28 multi_7x28_mod_5844(clk,rst,matrix_A[5844],matrix_B[44],mul_res1[5844]);
multi_7x28 multi_7x28_mod_5845(clk,rst,matrix_A[5845],matrix_B[45],mul_res1[5845]);
multi_7x28 multi_7x28_mod_5846(clk,rst,matrix_A[5846],matrix_B[46],mul_res1[5846]);
multi_7x28 multi_7x28_mod_5847(clk,rst,matrix_A[5847],matrix_B[47],mul_res1[5847]);
multi_7x28 multi_7x28_mod_5848(clk,rst,matrix_A[5848],matrix_B[48],mul_res1[5848]);
multi_7x28 multi_7x28_mod_5849(clk,rst,matrix_A[5849],matrix_B[49],mul_res1[5849]);
multi_7x28 multi_7x28_mod_5850(clk,rst,matrix_A[5850],matrix_B[50],mul_res1[5850]);
multi_7x28 multi_7x28_mod_5851(clk,rst,matrix_A[5851],matrix_B[51],mul_res1[5851]);
multi_7x28 multi_7x28_mod_5852(clk,rst,matrix_A[5852],matrix_B[52],mul_res1[5852]);
multi_7x28 multi_7x28_mod_5853(clk,rst,matrix_A[5853],matrix_B[53],mul_res1[5853]);
multi_7x28 multi_7x28_mod_5854(clk,rst,matrix_A[5854],matrix_B[54],mul_res1[5854]);
multi_7x28 multi_7x28_mod_5855(clk,rst,matrix_A[5855],matrix_B[55],mul_res1[5855]);
multi_7x28 multi_7x28_mod_5856(clk,rst,matrix_A[5856],matrix_B[56],mul_res1[5856]);
multi_7x28 multi_7x28_mod_5857(clk,rst,matrix_A[5857],matrix_B[57],mul_res1[5857]);
multi_7x28 multi_7x28_mod_5858(clk,rst,matrix_A[5858],matrix_B[58],mul_res1[5858]);
multi_7x28 multi_7x28_mod_5859(clk,rst,matrix_A[5859],matrix_B[59],mul_res1[5859]);
multi_7x28 multi_7x28_mod_5860(clk,rst,matrix_A[5860],matrix_B[60],mul_res1[5860]);
multi_7x28 multi_7x28_mod_5861(clk,rst,matrix_A[5861],matrix_B[61],mul_res1[5861]);
multi_7x28 multi_7x28_mod_5862(clk,rst,matrix_A[5862],matrix_B[62],mul_res1[5862]);
multi_7x28 multi_7x28_mod_5863(clk,rst,matrix_A[5863],matrix_B[63],mul_res1[5863]);
multi_7x28 multi_7x28_mod_5864(clk,rst,matrix_A[5864],matrix_B[64],mul_res1[5864]);
multi_7x28 multi_7x28_mod_5865(clk,rst,matrix_A[5865],matrix_B[65],mul_res1[5865]);
multi_7x28 multi_7x28_mod_5866(clk,rst,matrix_A[5866],matrix_B[66],mul_res1[5866]);
multi_7x28 multi_7x28_mod_5867(clk,rst,matrix_A[5867],matrix_B[67],mul_res1[5867]);
multi_7x28 multi_7x28_mod_5868(clk,rst,matrix_A[5868],matrix_B[68],mul_res1[5868]);
multi_7x28 multi_7x28_mod_5869(clk,rst,matrix_A[5869],matrix_B[69],mul_res1[5869]);
multi_7x28 multi_7x28_mod_5870(clk,rst,matrix_A[5870],matrix_B[70],mul_res1[5870]);
multi_7x28 multi_7x28_mod_5871(clk,rst,matrix_A[5871],matrix_B[71],mul_res1[5871]);
multi_7x28 multi_7x28_mod_5872(clk,rst,matrix_A[5872],matrix_B[72],mul_res1[5872]);
multi_7x28 multi_7x28_mod_5873(clk,rst,matrix_A[5873],matrix_B[73],mul_res1[5873]);
multi_7x28 multi_7x28_mod_5874(clk,rst,matrix_A[5874],matrix_B[74],mul_res1[5874]);
multi_7x28 multi_7x28_mod_5875(clk,rst,matrix_A[5875],matrix_B[75],mul_res1[5875]);
multi_7x28 multi_7x28_mod_5876(clk,rst,matrix_A[5876],matrix_B[76],mul_res1[5876]);
multi_7x28 multi_7x28_mod_5877(clk,rst,matrix_A[5877],matrix_B[77],mul_res1[5877]);
multi_7x28 multi_7x28_mod_5878(clk,rst,matrix_A[5878],matrix_B[78],mul_res1[5878]);
multi_7x28 multi_7x28_mod_5879(clk,rst,matrix_A[5879],matrix_B[79],mul_res1[5879]);
multi_7x28 multi_7x28_mod_5880(clk,rst,matrix_A[5880],matrix_B[80],mul_res1[5880]);
multi_7x28 multi_7x28_mod_5881(clk,rst,matrix_A[5881],matrix_B[81],mul_res1[5881]);
multi_7x28 multi_7x28_mod_5882(clk,rst,matrix_A[5882],matrix_B[82],mul_res1[5882]);
multi_7x28 multi_7x28_mod_5883(clk,rst,matrix_A[5883],matrix_B[83],mul_res1[5883]);
multi_7x28 multi_7x28_mod_5884(clk,rst,matrix_A[5884],matrix_B[84],mul_res1[5884]);
multi_7x28 multi_7x28_mod_5885(clk,rst,matrix_A[5885],matrix_B[85],mul_res1[5885]);
multi_7x28 multi_7x28_mod_5886(clk,rst,matrix_A[5886],matrix_B[86],mul_res1[5886]);
multi_7x28 multi_7x28_mod_5887(clk,rst,matrix_A[5887],matrix_B[87],mul_res1[5887]);
multi_7x28 multi_7x28_mod_5888(clk,rst,matrix_A[5888],matrix_B[88],mul_res1[5888]);
multi_7x28 multi_7x28_mod_5889(clk,rst,matrix_A[5889],matrix_B[89],mul_res1[5889]);
multi_7x28 multi_7x28_mod_5890(clk,rst,matrix_A[5890],matrix_B[90],mul_res1[5890]);
multi_7x28 multi_7x28_mod_5891(clk,rst,matrix_A[5891],matrix_B[91],mul_res1[5891]);
multi_7x28 multi_7x28_mod_5892(clk,rst,matrix_A[5892],matrix_B[92],mul_res1[5892]);
multi_7x28 multi_7x28_mod_5893(clk,rst,matrix_A[5893],matrix_B[93],mul_res1[5893]);
multi_7x28 multi_7x28_mod_5894(clk,rst,matrix_A[5894],matrix_B[94],mul_res1[5894]);
multi_7x28 multi_7x28_mod_5895(clk,rst,matrix_A[5895],matrix_B[95],mul_res1[5895]);
multi_7x28 multi_7x28_mod_5896(clk,rst,matrix_A[5896],matrix_B[96],mul_res1[5896]);
multi_7x28 multi_7x28_mod_5897(clk,rst,matrix_A[5897],matrix_B[97],mul_res1[5897]);
multi_7x28 multi_7x28_mod_5898(clk,rst,matrix_A[5898],matrix_B[98],mul_res1[5898]);
multi_7x28 multi_7x28_mod_5899(clk,rst,matrix_A[5899],matrix_B[99],mul_res1[5899]);
multi_7x28 multi_7x28_mod_5900(clk,rst,matrix_A[5900],matrix_B[100],mul_res1[5900]);
multi_7x28 multi_7x28_mod_5901(clk,rst,matrix_A[5901],matrix_B[101],mul_res1[5901]);
multi_7x28 multi_7x28_mod_5902(clk,rst,matrix_A[5902],matrix_B[102],mul_res1[5902]);
multi_7x28 multi_7x28_mod_5903(clk,rst,matrix_A[5903],matrix_B[103],mul_res1[5903]);
multi_7x28 multi_7x28_mod_5904(clk,rst,matrix_A[5904],matrix_B[104],mul_res1[5904]);
multi_7x28 multi_7x28_mod_5905(clk,rst,matrix_A[5905],matrix_B[105],mul_res1[5905]);
multi_7x28 multi_7x28_mod_5906(clk,rst,matrix_A[5906],matrix_B[106],mul_res1[5906]);
multi_7x28 multi_7x28_mod_5907(clk,rst,matrix_A[5907],matrix_B[107],mul_res1[5907]);
multi_7x28 multi_7x28_mod_5908(clk,rst,matrix_A[5908],matrix_B[108],mul_res1[5908]);
multi_7x28 multi_7x28_mod_5909(clk,rst,matrix_A[5909],matrix_B[109],mul_res1[5909]);
multi_7x28 multi_7x28_mod_5910(clk,rst,matrix_A[5910],matrix_B[110],mul_res1[5910]);
multi_7x28 multi_7x28_mod_5911(clk,rst,matrix_A[5911],matrix_B[111],mul_res1[5911]);
multi_7x28 multi_7x28_mod_5912(clk,rst,matrix_A[5912],matrix_B[112],mul_res1[5912]);
multi_7x28 multi_7x28_mod_5913(clk,rst,matrix_A[5913],matrix_B[113],mul_res1[5913]);
multi_7x28 multi_7x28_mod_5914(clk,rst,matrix_A[5914],matrix_B[114],mul_res1[5914]);
multi_7x28 multi_7x28_mod_5915(clk,rst,matrix_A[5915],matrix_B[115],mul_res1[5915]);
multi_7x28 multi_7x28_mod_5916(clk,rst,matrix_A[5916],matrix_B[116],mul_res1[5916]);
multi_7x28 multi_7x28_mod_5917(clk,rst,matrix_A[5917],matrix_B[117],mul_res1[5917]);
multi_7x28 multi_7x28_mod_5918(clk,rst,matrix_A[5918],matrix_B[118],mul_res1[5918]);
multi_7x28 multi_7x28_mod_5919(clk,rst,matrix_A[5919],matrix_B[119],mul_res1[5919]);
multi_7x28 multi_7x28_mod_5920(clk,rst,matrix_A[5920],matrix_B[120],mul_res1[5920]);
multi_7x28 multi_7x28_mod_5921(clk,rst,matrix_A[5921],matrix_B[121],mul_res1[5921]);
multi_7x28 multi_7x28_mod_5922(clk,rst,matrix_A[5922],matrix_B[122],mul_res1[5922]);
multi_7x28 multi_7x28_mod_5923(clk,rst,matrix_A[5923],matrix_B[123],mul_res1[5923]);
multi_7x28 multi_7x28_mod_5924(clk,rst,matrix_A[5924],matrix_B[124],mul_res1[5924]);
multi_7x28 multi_7x28_mod_5925(clk,rst,matrix_A[5925],matrix_B[125],mul_res1[5925]);
multi_7x28 multi_7x28_mod_5926(clk,rst,matrix_A[5926],matrix_B[126],mul_res1[5926]);
multi_7x28 multi_7x28_mod_5927(clk,rst,matrix_A[5927],matrix_B[127],mul_res1[5927]);
multi_7x28 multi_7x28_mod_5928(clk,rst,matrix_A[5928],matrix_B[128],mul_res1[5928]);
multi_7x28 multi_7x28_mod_5929(clk,rst,matrix_A[5929],matrix_B[129],mul_res1[5929]);
multi_7x28 multi_7x28_mod_5930(clk,rst,matrix_A[5930],matrix_B[130],mul_res1[5930]);
multi_7x28 multi_7x28_mod_5931(clk,rst,matrix_A[5931],matrix_B[131],mul_res1[5931]);
multi_7x28 multi_7x28_mod_5932(clk,rst,matrix_A[5932],matrix_B[132],mul_res1[5932]);
multi_7x28 multi_7x28_mod_5933(clk,rst,matrix_A[5933],matrix_B[133],mul_res1[5933]);
multi_7x28 multi_7x28_mod_5934(clk,rst,matrix_A[5934],matrix_B[134],mul_res1[5934]);
multi_7x28 multi_7x28_mod_5935(clk,rst,matrix_A[5935],matrix_B[135],mul_res1[5935]);
multi_7x28 multi_7x28_mod_5936(clk,rst,matrix_A[5936],matrix_B[136],mul_res1[5936]);
multi_7x28 multi_7x28_mod_5937(clk,rst,matrix_A[5937],matrix_B[137],mul_res1[5937]);
multi_7x28 multi_7x28_mod_5938(clk,rst,matrix_A[5938],matrix_B[138],mul_res1[5938]);
multi_7x28 multi_7x28_mod_5939(clk,rst,matrix_A[5939],matrix_B[139],mul_res1[5939]);
multi_7x28 multi_7x28_mod_5940(clk,rst,matrix_A[5940],matrix_B[140],mul_res1[5940]);
multi_7x28 multi_7x28_mod_5941(clk,rst,matrix_A[5941],matrix_B[141],mul_res1[5941]);
multi_7x28 multi_7x28_mod_5942(clk,rst,matrix_A[5942],matrix_B[142],mul_res1[5942]);
multi_7x28 multi_7x28_mod_5943(clk,rst,matrix_A[5943],matrix_B[143],mul_res1[5943]);
multi_7x28 multi_7x28_mod_5944(clk,rst,matrix_A[5944],matrix_B[144],mul_res1[5944]);
multi_7x28 multi_7x28_mod_5945(clk,rst,matrix_A[5945],matrix_B[145],mul_res1[5945]);
multi_7x28 multi_7x28_mod_5946(clk,rst,matrix_A[5946],matrix_B[146],mul_res1[5946]);
multi_7x28 multi_7x28_mod_5947(clk,rst,matrix_A[5947],matrix_B[147],mul_res1[5947]);
multi_7x28 multi_7x28_mod_5948(clk,rst,matrix_A[5948],matrix_B[148],mul_res1[5948]);
multi_7x28 multi_7x28_mod_5949(clk,rst,matrix_A[5949],matrix_B[149],mul_res1[5949]);
multi_7x28 multi_7x28_mod_5950(clk,rst,matrix_A[5950],matrix_B[150],mul_res1[5950]);
multi_7x28 multi_7x28_mod_5951(clk,rst,matrix_A[5951],matrix_B[151],mul_res1[5951]);
multi_7x28 multi_7x28_mod_5952(clk,rst,matrix_A[5952],matrix_B[152],mul_res1[5952]);
multi_7x28 multi_7x28_mod_5953(clk,rst,matrix_A[5953],matrix_B[153],mul_res1[5953]);
multi_7x28 multi_7x28_mod_5954(clk,rst,matrix_A[5954],matrix_B[154],mul_res1[5954]);
multi_7x28 multi_7x28_mod_5955(clk,rst,matrix_A[5955],matrix_B[155],mul_res1[5955]);
multi_7x28 multi_7x28_mod_5956(clk,rst,matrix_A[5956],matrix_B[156],mul_res1[5956]);
multi_7x28 multi_7x28_mod_5957(clk,rst,matrix_A[5957],matrix_B[157],mul_res1[5957]);
multi_7x28 multi_7x28_mod_5958(clk,rst,matrix_A[5958],matrix_B[158],mul_res1[5958]);
multi_7x28 multi_7x28_mod_5959(clk,rst,matrix_A[5959],matrix_B[159],mul_res1[5959]);
multi_7x28 multi_7x28_mod_5960(clk,rst,matrix_A[5960],matrix_B[160],mul_res1[5960]);
multi_7x28 multi_7x28_mod_5961(clk,rst,matrix_A[5961],matrix_B[161],mul_res1[5961]);
multi_7x28 multi_7x28_mod_5962(clk,rst,matrix_A[5962],matrix_B[162],mul_res1[5962]);
multi_7x28 multi_7x28_mod_5963(clk,rst,matrix_A[5963],matrix_B[163],mul_res1[5963]);
multi_7x28 multi_7x28_mod_5964(clk,rst,matrix_A[5964],matrix_B[164],mul_res1[5964]);
multi_7x28 multi_7x28_mod_5965(clk,rst,matrix_A[5965],matrix_B[165],mul_res1[5965]);
multi_7x28 multi_7x28_mod_5966(clk,rst,matrix_A[5966],matrix_B[166],mul_res1[5966]);
multi_7x28 multi_7x28_mod_5967(clk,rst,matrix_A[5967],matrix_B[167],mul_res1[5967]);
multi_7x28 multi_7x28_mod_5968(clk,rst,matrix_A[5968],matrix_B[168],mul_res1[5968]);
multi_7x28 multi_7x28_mod_5969(clk,rst,matrix_A[5969],matrix_B[169],mul_res1[5969]);
multi_7x28 multi_7x28_mod_5970(clk,rst,matrix_A[5970],matrix_B[170],mul_res1[5970]);
multi_7x28 multi_7x28_mod_5971(clk,rst,matrix_A[5971],matrix_B[171],mul_res1[5971]);
multi_7x28 multi_7x28_mod_5972(clk,rst,matrix_A[5972],matrix_B[172],mul_res1[5972]);
multi_7x28 multi_7x28_mod_5973(clk,rst,matrix_A[5973],matrix_B[173],mul_res1[5973]);
multi_7x28 multi_7x28_mod_5974(clk,rst,matrix_A[5974],matrix_B[174],mul_res1[5974]);
multi_7x28 multi_7x28_mod_5975(clk,rst,matrix_A[5975],matrix_B[175],mul_res1[5975]);
multi_7x28 multi_7x28_mod_5976(clk,rst,matrix_A[5976],matrix_B[176],mul_res1[5976]);
multi_7x28 multi_7x28_mod_5977(clk,rst,matrix_A[5977],matrix_B[177],mul_res1[5977]);
multi_7x28 multi_7x28_mod_5978(clk,rst,matrix_A[5978],matrix_B[178],mul_res1[5978]);
multi_7x28 multi_7x28_mod_5979(clk,rst,matrix_A[5979],matrix_B[179],mul_res1[5979]);
multi_7x28 multi_7x28_mod_5980(clk,rst,matrix_A[5980],matrix_B[180],mul_res1[5980]);
multi_7x28 multi_7x28_mod_5981(clk,rst,matrix_A[5981],matrix_B[181],mul_res1[5981]);
multi_7x28 multi_7x28_mod_5982(clk,rst,matrix_A[5982],matrix_B[182],mul_res1[5982]);
multi_7x28 multi_7x28_mod_5983(clk,rst,matrix_A[5983],matrix_B[183],mul_res1[5983]);
multi_7x28 multi_7x28_mod_5984(clk,rst,matrix_A[5984],matrix_B[184],mul_res1[5984]);
multi_7x28 multi_7x28_mod_5985(clk,rst,matrix_A[5985],matrix_B[185],mul_res1[5985]);
multi_7x28 multi_7x28_mod_5986(clk,rst,matrix_A[5986],matrix_B[186],mul_res1[5986]);
multi_7x28 multi_7x28_mod_5987(clk,rst,matrix_A[5987],matrix_B[187],mul_res1[5987]);
multi_7x28 multi_7x28_mod_5988(clk,rst,matrix_A[5988],matrix_B[188],mul_res1[5988]);
multi_7x28 multi_7x28_mod_5989(clk,rst,matrix_A[5989],matrix_B[189],mul_res1[5989]);
multi_7x28 multi_7x28_mod_5990(clk,rst,matrix_A[5990],matrix_B[190],mul_res1[5990]);
multi_7x28 multi_7x28_mod_5991(clk,rst,matrix_A[5991],matrix_B[191],mul_res1[5991]);
multi_7x28 multi_7x28_mod_5992(clk,rst,matrix_A[5992],matrix_B[192],mul_res1[5992]);
multi_7x28 multi_7x28_mod_5993(clk,rst,matrix_A[5993],matrix_B[193],mul_res1[5993]);
multi_7x28 multi_7x28_mod_5994(clk,rst,matrix_A[5994],matrix_B[194],mul_res1[5994]);
multi_7x28 multi_7x28_mod_5995(clk,rst,matrix_A[5995],matrix_B[195],mul_res1[5995]);
multi_7x28 multi_7x28_mod_5996(clk,rst,matrix_A[5996],matrix_B[196],mul_res1[5996]);
multi_7x28 multi_7x28_mod_5997(clk,rst,matrix_A[5997],matrix_B[197],mul_res1[5997]);
multi_7x28 multi_7x28_mod_5998(clk,rst,matrix_A[5998],matrix_B[198],mul_res1[5998]);
multi_7x28 multi_7x28_mod_5999(clk,rst,matrix_A[5999],matrix_B[199],mul_res1[5999]);
multi_7x28 multi_7x28_mod_6000(clk,rst,matrix_A[6000],matrix_B[0],mul_res1[6000]);
multi_7x28 multi_7x28_mod_6001(clk,rst,matrix_A[6001],matrix_B[1],mul_res1[6001]);
multi_7x28 multi_7x28_mod_6002(clk,rst,matrix_A[6002],matrix_B[2],mul_res1[6002]);
multi_7x28 multi_7x28_mod_6003(clk,rst,matrix_A[6003],matrix_B[3],mul_res1[6003]);
multi_7x28 multi_7x28_mod_6004(clk,rst,matrix_A[6004],matrix_B[4],mul_res1[6004]);
multi_7x28 multi_7x28_mod_6005(clk,rst,matrix_A[6005],matrix_B[5],mul_res1[6005]);
multi_7x28 multi_7x28_mod_6006(clk,rst,matrix_A[6006],matrix_B[6],mul_res1[6006]);
multi_7x28 multi_7x28_mod_6007(clk,rst,matrix_A[6007],matrix_B[7],mul_res1[6007]);
multi_7x28 multi_7x28_mod_6008(clk,rst,matrix_A[6008],matrix_B[8],mul_res1[6008]);
multi_7x28 multi_7x28_mod_6009(clk,rst,matrix_A[6009],matrix_B[9],mul_res1[6009]);
multi_7x28 multi_7x28_mod_6010(clk,rst,matrix_A[6010],matrix_B[10],mul_res1[6010]);
multi_7x28 multi_7x28_mod_6011(clk,rst,matrix_A[6011],matrix_B[11],mul_res1[6011]);
multi_7x28 multi_7x28_mod_6012(clk,rst,matrix_A[6012],matrix_B[12],mul_res1[6012]);
multi_7x28 multi_7x28_mod_6013(clk,rst,matrix_A[6013],matrix_B[13],mul_res1[6013]);
multi_7x28 multi_7x28_mod_6014(clk,rst,matrix_A[6014],matrix_B[14],mul_res1[6014]);
multi_7x28 multi_7x28_mod_6015(clk,rst,matrix_A[6015],matrix_B[15],mul_res1[6015]);
multi_7x28 multi_7x28_mod_6016(clk,rst,matrix_A[6016],matrix_B[16],mul_res1[6016]);
multi_7x28 multi_7x28_mod_6017(clk,rst,matrix_A[6017],matrix_B[17],mul_res1[6017]);
multi_7x28 multi_7x28_mod_6018(clk,rst,matrix_A[6018],matrix_B[18],mul_res1[6018]);
multi_7x28 multi_7x28_mod_6019(clk,rst,matrix_A[6019],matrix_B[19],mul_res1[6019]);
multi_7x28 multi_7x28_mod_6020(clk,rst,matrix_A[6020],matrix_B[20],mul_res1[6020]);
multi_7x28 multi_7x28_mod_6021(clk,rst,matrix_A[6021],matrix_B[21],mul_res1[6021]);
multi_7x28 multi_7x28_mod_6022(clk,rst,matrix_A[6022],matrix_B[22],mul_res1[6022]);
multi_7x28 multi_7x28_mod_6023(clk,rst,matrix_A[6023],matrix_B[23],mul_res1[6023]);
multi_7x28 multi_7x28_mod_6024(clk,rst,matrix_A[6024],matrix_B[24],mul_res1[6024]);
multi_7x28 multi_7x28_mod_6025(clk,rst,matrix_A[6025],matrix_B[25],mul_res1[6025]);
multi_7x28 multi_7x28_mod_6026(clk,rst,matrix_A[6026],matrix_B[26],mul_res1[6026]);
multi_7x28 multi_7x28_mod_6027(clk,rst,matrix_A[6027],matrix_B[27],mul_res1[6027]);
multi_7x28 multi_7x28_mod_6028(clk,rst,matrix_A[6028],matrix_B[28],mul_res1[6028]);
multi_7x28 multi_7x28_mod_6029(clk,rst,matrix_A[6029],matrix_B[29],mul_res1[6029]);
multi_7x28 multi_7x28_mod_6030(clk,rst,matrix_A[6030],matrix_B[30],mul_res1[6030]);
multi_7x28 multi_7x28_mod_6031(clk,rst,matrix_A[6031],matrix_B[31],mul_res1[6031]);
multi_7x28 multi_7x28_mod_6032(clk,rst,matrix_A[6032],matrix_B[32],mul_res1[6032]);
multi_7x28 multi_7x28_mod_6033(clk,rst,matrix_A[6033],matrix_B[33],mul_res1[6033]);
multi_7x28 multi_7x28_mod_6034(clk,rst,matrix_A[6034],matrix_B[34],mul_res1[6034]);
multi_7x28 multi_7x28_mod_6035(clk,rst,matrix_A[6035],matrix_B[35],mul_res1[6035]);
multi_7x28 multi_7x28_mod_6036(clk,rst,matrix_A[6036],matrix_B[36],mul_res1[6036]);
multi_7x28 multi_7x28_mod_6037(clk,rst,matrix_A[6037],matrix_B[37],mul_res1[6037]);
multi_7x28 multi_7x28_mod_6038(clk,rst,matrix_A[6038],matrix_B[38],mul_res1[6038]);
multi_7x28 multi_7x28_mod_6039(clk,rst,matrix_A[6039],matrix_B[39],mul_res1[6039]);
multi_7x28 multi_7x28_mod_6040(clk,rst,matrix_A[6040],matrix_B[40],mul_res1[6040]);
multi_7x28 multi_7x28_mod_6041(clk,rst,matrix_A[6041],matrix_B[41],mul_res1[6041]);
multi_7x28 multi_7x28_mod_6042(clk,rst,matrix_A[6042],matrix_B[42],mul_res1[6042]);
multi_7x28 multi_7x28_mod_6043(clk,rst,matrix_A[6043],matrix_B[43],mul_res1[6043]);
multi_7x28 multi_7x28_mod_6044(clk,rst,matrix_A[6044],matrix_B[44],mul_res1[6044]);
multi_7x28 multi_7x28_mod_6045(clk,rst,matrix_A[6045],matrix_B[45],mul_res1[6045]);
multi_7x28 multi_7x28_mod_6046(clk,rst,matrix_A[6046],matrix_B[46],mul_res1[6046]);
multi_7x28 multi_7x28_mod_6047(clk,rst,matrix_A[6047],matrix_B[47],mul_res1[6047]);
multi_7x28 multi_7x28_mod_6048(clk,rst,matrix_A[6048],matrix_B[48],mul_res1[6048]);
multi_7x28 multi_7x28_mod_6049(clk,rst,matrix_A[6049],matrix_B[49],mul_res1[6049]);
multi_7x28 multi_7x28_mod_6050(clk,rst,matrix_A[6050],matrix_B[50],mul_res1[6050]);
multi_7x28 multi_7x28_mod_6051(clk,rst,matrix_A[6051],matrix_B[51],mul_res1[6051]);
multi_7x28 multi_7x28_mod_6052(clk,rst,matrix_A[6052],matrix_B[52],mul_res1[6052]);
multi_7x28 multi_7x28_mod_6053(clk,rst,matrix_A[6053],matrix_B[53],mul_res1[6053]);
multi_7x28 multi_7x28_mod_6054(clk,rst,matrix_A[6054],matrix_B[54],mul_res1[6054]);
multi_7x28 multi_7x28_mod_6055(clk,rst,matrix_A[6055],matrix_B[55],mul_res1[6055]);
multi_7x28 multi_7x28_mod_6056(clk,rst,matrix_A[6056],matrix_B[56],mul_res1[6056]);
multi_7x28 multi_7x28_mod_6057(clk,rst,matrix_A[6057],matrix_B[57],mul_res1[6057]);
multi_7x28 multi_7x28_mod_6058(clk,rst,matrix_A[6058],matrix_B[58],mul_res1[6058]);
multi_7x28 multi_7x28_mod_6059(clk,rst,matrix_A[6059],matrix_B[59],mul_res1[6059]);
multi_7x28 multi_7x28_mod_6060(clk,rst,matrix_A[6060],matrix_B[60],mul_res1[6060]);
multi_7x28 multi_7x28_mod_6061(clk,rst,matrix_A[6061],matrix_B[61],mul_res1[6061]);
multi_7x28 multi_7x28_mod_6062(clk,rst,matrix_A[6062],matrix_B[62],mul_res1[6062]);
multi_7x28 multi_7x28_mod_6063(clk,rst,matrix_A[6063],matrix_B[63],mul_res1[6063]);
multi_7x28 multi_7x28_mod_6064(clk,rst,matrix_A[6064],matrix_B[64],mul_res1[6064]);
multi_7x28 multi_7x28_mod_6065(clk,rst,matrix_A[6065],matrix_B[65],mul_res1[6065]);
multi_7x28 multi_7x28_mod_6066(clk,rst,matrix_A[6066],matrix_B[66],mul_res1[6066]);
multi_7x28 multi_7x28_mod_6067(clk,rst,matrix_A[6067],matrix_B[67],mul_res1[6067]);
multi_7x28 multi_7x28_mod_6068(clk,rst,matrix_A[6068],matrix_B[68],mul_res1[6068]);
multi_7x28 multi_7x28_mod_6069(clk,rst,matrix_A[6069],matrix_B[69],mul_res1[6069]);
multi_7x28 multi_7x28_mod_6070(clk,rst,matrix_A[6070],matrix_B[70],mul_res1[6070]);
multi_7x28 multi_7x28_mod_6071(clk,rst,matrix_A[6071],matrix_B[71],mul_res1[6071]);
multi_7x28 multi_7x28_mod_6072(clk,rst,matrix_A[6072],matrix_B[72],mul_res1[6072]);
multi_7x28 multi_7x28_mod_6073(clk,rst,matrix_A[6073],matrix_B[73],mul_res1[6073]);
multi_7x28 multi_7x28_mod_6074(clk,rst,matrix_A[6074],matrix_B[74],mul_res1[6074]);
multi_7x28 multi_7x28_mod_6075(clk,rst,matrix_A[6075],matrix_B[75],mul_res1[6075]);
multi_7x28 multi_7x28_mod_6076(clk,rst,matrix_A[6076],matrix_B[76],mul_res1[6076]);
multi_7x28 multi_7x28_mod_6077(clk,rst,matrix_A[6077],matrix_B[77],mul_res1[6077]);
multi_7x28 multi_7x28_mod_6078(clk,rst,matrix_A[6078],matrix_B[78],mul_res1[6078]);
multi_7x28 multi_7x28_mod_6079(clk,rst,matrix_A[6079],matrix_B[79],mul_res1[6079]);
multi_7x28 multi_7x28_mod_6080(clk,rst,matrix_A[6080],matrix_B[80],mul_res1[6080]);
multi_7x28 multi_7x28_mod_6081(clk,rst,matrix_A[6081],matrix_B[81],mul_res1[6081]);
multi_7x28 multi_7x28_mod_6082(clk,rst,matrix_A[6082],matrix_B[82],mul_res1[6082]);
multi_7x28 multi_7x28_mod_6083(clk,rst,matrix_A[6083],matrix_B[83],mul_res1[6083]);
multi_7x28 multi_7x28_mod_6084(clk,rst,matrix_A[6084],matrix_B[84],mul_res1[6084]);
multi_7x28 multi_7x28_mod_6085(clk,rst,matrix_A[6085],matrix_B[85],mul_res1[6085]);
multi_7x28 multi_7x28_mod_6086(clk,rst,matrix_A[6086],matrix_B[86],mul_res1[6086]);
multi_7x28 multi_7x28_mod_6087(clk,rst,matrix_A[6087],matrix_B[87],mul_res1[6087]);
multi_7x28 multi_7x28_mod_6088(clk,rst,matrix_A[6088],matrix_B[88],mul_res1[6088]);
multi_7x28 multi_7x28_mod_6089(clk,rst,matrix_A[6089],matrix_B[89],mul_res1[6089]);
multi_7x28 multi_7x28_mod_6090(clk,rst,matrix_A[6090],matrix_B[90],mul_res1[6090]);
multi_7x28 multi_7x28_mod_6091(clk,rst,matrix_A[6091],matrix_B[91],mul_res1[6091]);
multi_7x28 multi_7x28_mod_6092(clk,rst,matrix_A[6092],matrix_B[92],mul_res1[6092]);
multi_7x28 multi_7x28_mod_6093(clk,rst,matrix_A[6093],matrix_B[93],mul_res1[6093]);
multi_7x28 multi_7x28_mod_6094(clk,rst,matrix_A[6094],matrix_B[94],mul_res1[6094]);
multi_7x28 multi_7x28_mod_6095(clk,rst,matrix_A[6095],matrix_B[95],mul_res1[6095]);
multi_7x28 multi_7x28_mod_6096(clk,rst,matrix_A[6096],matrix_B[96],mul_res1[6096]);
multi_7x28 multi_7x28_mod_6097(clk,rst,matrix_A[6097],matrix_B[97],mul_res1[6097]);
multi_7x28 multi_7x28_mod_6098(clk,rst,matrix_A[6098],matrix_B[98],mul_res1[6098]);
multi_7x28 multi_7x28_mod_6099(clk,rst,matrix_A[6099],matrix_B[99],mul_res1[6099]);
multi_7x28 multi_7x28_mod_6100(clk,rst,matrix_A[6100],matrix_B[100],mul_res1[6100]);
multi_7x28 multi_7x28_mod_6101(clk,rst,matrix_A[6101],matrix_B[101],mul_res1[6101]);
multi_7x28 multi_7x28_mod_6102(clk,rst,matrix_A[6102],matrix_B[102],mul_res1[6102]);
multi_7x28 multi_7x28_mod_6103(clk,rst,matrix_A[6103],matrix_B[103],mul_res1[6103]);
multi_7x28 multi_7x28_mod_6104(clk,rst,matrix_A[6104],matrix_B[104],mul_res1[6104]);
multi_7x28 multi_7x28_mod_6105(clk,rst,matrix_A[6105],matrix_B[105],mul_res1[6105]);
multi_7x28 multi_7x28_mod_6106(clk,rst,matrix_A[6106],matrix_B[106],mul_res1[6106]);
multi_7x28 multi_7x28_mod_6107(clk,rst,matrix_A[6107],matrix_B[107],mul_res1[6107]);
multi_7x28 multi_7x28_mod_6108(clk,rst,matrix_A[6108],matrix_B[108],mul_res1[6108]);
multi_7x28 multi_7x28_mod_6109(clk,rst,matrix_A[6109],matrix_B[109],mul_res1[6109]);
multi_7x28 multi_7x28_mod_6110(clk,rst,matrix_A[6110],matrix_B[110],mul_res1[6110]);
multi_7x28 multi_7x28_mod_6111(clk,rst,matrix_A[6111],matrix_B[111],mul_res1[6111]);
multi_7x28 multi_7x28_mod_6112(clk,rst,matrix_A[6112],matrix_B[112],mul_res1[6112]);
multi_7x28 multi_7x28_mod_6113(clk,rst,matrix_A[6113],matrix_B[113],mul_res1[6113]);
multi_7x28 multi_7x28_mod_6114(clk,rst,matrix_A[6114],matrix_B[114],mul_res1[6114]);
multi_7x28 multi_7x28_mod_6115(clk,rst,matrix_A[6115],matrix_B[115],mul_res1[6115]);
multi_7x28 multi_7x28_mod_6116(clk,rst,matrix_A[6116],matrix_B[116],mul_res1[6116]);
multi_7x28 multi_7x28_mod_6117(clk,rst,matrix_A[6117],matrix_B[117],mul_res1[6117]);
multi_7x28 multi_7x28_mod_6118(clk,rst,matrix_A[6118],matrix_B[118],mul_res1[6118]);
multi_7x28 multi_7x28_mod_6119(clk,rst,matrix_A[6119],matrix_B[119],mul_res1[6119]);
multi_7x28 multi_7x28_mod_6120(clk,rst,matrix_A[6120],matrix_B[120],mul_res1[6120]);
multi_7x28 multi_7x28_mod_6121(clk,rst,matrix_A[6121],matrix_B[121],mul_res1[6121]);
multi_7x28 multi_7x28_mod_6122(clk,rst,matrix_A[6122],matrix_B[122],mul_res1[6122]);
multi_7x28 multi_7x28_mod_6123(clk,rst,matrix_A[6123],matrix_B[123],mul_res1[6123]);
multi_7x28 multi_7x28_mod_6124(clk,rst,matrix_A[6124],matrix_B[124],mul_res1[6124]);
multi_7x28 multi_7x28_mod_6125(clk,rst,matrix_A[6125],matrix_B[125],mul_res1[6125]);
multi_7x28 multi_7x28_mod_6126(clk,rst,matrix_A[6126],matrix_B[126],mul_res1[6126]);
multi_7x28 multi_7x28_mod_6127(clk,rst,matrix_A[6127],matrix_B[127],mul_res1[6127]);
multi_7x28 multi_7x28_mod_6128(clk,rst,matrix_A[6128],matrix_B[128],mul_res1[6128]);
multi_7x28 multi_7x28_mod_6129(clk,rst,matrix_A[6129],matrix_B[129],mul_res1[6129]);
multi_7x28 multi_7x28_mod_6130(clk,rst,matrix_A[6130],matrix_B[130],mul_res1[6130]);
multi_7x28 multi_7x28_mod_6131(clk,rst,matrix_A[6131],matrix_B[131],mul_res1[6131]);
multi_7x28 multi_7x28_mod_6132(clk,rst,matrix_A[6132],matrix_B[132],mul_res1[6132]);
multi_7x28 multi_7x28_mod_6133(clk,rst,matrix_A[6133],matrix_B[133],mul_res1[6133]);
multi_7x28 multi_7x28_mod_6134(clk,rst,matrix_A[6134],matrix_B[134],mul_res1[6134]);
multi_7x28 multi_7x28_mod_6135(clk,rst,matrix_A[6135],matrix_B[135],mul_res1[6135]);
multi_7x28 multi_7x28_mod_6136(clk,rst,matrix_A[6136],matrix_B[136],mul_res1[6136]);
multi_7x28 multi_7x28_mod_6137(clk,rst,matrix_A[6137],matrix_B[137],mul_res1[6137]);
multi_7x28 multi_7x28_mod_6138(clk,rst,matrix_A[6138],matrix_B[138],mul_res1[6138]);
multi_7x28 multi_7x28_mod_6139(clk,rst,matrix_A[6139],matrix_B[139],mul_res1[6139]);
multi_7x28 multi_7x28_mod_6140(clk,rst,matrix_A[6140],matrix_B[140],mul_res1[6140]);
multi_7x28 multi_7x28_mod_6141(clk,rst,matrix_A[6141],matrix_B[141],mul_res1[6141]);
multi_7x28 multi_7x28_mod_6142(clk,rst,matrix_A[6142],matrix_B[142],mul_res1[6142]);
multi_7x28 multi_7x28_mod_6143(clk,rst,matrix_A[6143],matrix_B[143],mul_res1[6143]);
multi_7x28 multi_7x28_mod_6144(clk,rst,matrix_A[6144],matrix_B[144],mul_res1[6144]);
multi_7x28 multi_7x28_mod_6145(clk,rst,matrix_A[6145],matrix_B[145],mul_res1[6145]);
multi_7x28 multi_7x28_mod_6146(clk,rst,matrix_A[6146],matrix_B[146],mul_res1[6146]);
multi_7x28 multi_7x28_mod_6147(clk,rst,matrix_A[6147],matrix_B[147],mul_res1[6147]);
multi_7x28 multi_7x28_mod_6148(clk,rst,matrix_A[6148],matrix_B[148],mul_res1[6148]);
multi_7x28 multi_7x28_mod_6149(clk,rst,matrix_A[6149],matrix_B[149],mul_res1[6149]);
multi_7x28 multi_7x28_mod_6150(clk,rst,matrix_A[6150],matrix_B[150],mul_res1[6150]);
multi_7x28 multi_7x28_mod_6151(clk,rst,matrix_A[6151],matrix_B[151],mul_res1[6151]);
multi_7x28 multi_7x28_mod_6152(clk,rst,matrix_A[6152],matrix_B[152],mul_res1[6152]);
multi_7x28 multi_7x28_mod_6153(clk,rst,matrix_A[6153],matrix_B[153],mul_res1[6153]);
multi_7x28 multi_7x28_mod_6154(clk,rst,matrix_A[6154],matrix_B[154],mul_res1[6154]);
multi_7x28 multi_7x28_mod_6155(clk,rst,matrix_A[6155],matrix_B[155],mul_res1[6155]);
multi_7x28 multi_7x28_mod_6156(clk,rst,matrix_A[6156],matrix_B[156],mul_res1[6156]);
multi_7x28 multi_7x28_mod_6157(clk,rst,matrix_A[6157],matrix_B[157],mul_res1[6157]);
multi_7x28 multi_7x28_mod_6158(clk,rst,matrix_A[6158],matrix_B[158],mul_res1[6158]);
multi_7x28 multi_7x28_mod_6159(clk,rst,matrix_A[6159],matrix_B[159],mul_res1[6159]);
multi_7x28 multi_7x28_mod_6160(clk,rst,matrix_A[6160],matrix_B[160],mul_res1[6160]);
multi_7x28 multi_7x28_mod_6161(clk,rst,matrix_A[6161],matrix_B[161],mul_res1[6161]);
multi_7x28 multi_7x28_mod_6162(clk,rst,matrix_A[6162],matrix_B[162],mul_res1[6162]);
multi_7x28 multi_7x28_mod_6163(clk,rst,matrix_A[6163],matrix_B[163],mul_res1[6163]);
multi_7x28 multi_7x28_mod_6164(clk,rst,matrix_A[6164],matrix_B[164],mul_res1[6164]);
multi_7x28 multi_7x28_mod_6165(clk,rst,matrix_A[6165],matrix_B[165],mul_res1[6165]);
multi_7x28 multi_7x28_mod_6166(clk,rst,matrix_A[6166],matrix_B[166],mul_res1[6166]);
multi_7x28 multi_7x28_mod_6167(clk,rst,matrix_A[6167],matrix_B[167],mul_res1[6167]);
multi_7x28 multi_7x28_mod_6168(clk,rst,matrix_A[6168],matrix_B[168],mul_res1[6168]);
multi_7x28 multi_7x28_mod_6169(clk,rst,matrix_A[6169],matrix_B[169],mul_res1[6169]);
multi_7x28 multi_7x28_mod_6170(clk,rst,matrix_A[6170],matrix_B[170],mul_res1[6170]);
multi_7x28 multi_7x28_mod_6171(clk,rst,matrix_A[6171],matrix_B[171],mul_res1[6171]);
multi_7x28 multi_7x28_mod_6172(clk,rst,matrix_A[6172],matrix_B[172],mul_res1[6172]);
multi_7x28 multi_7x28_mod_6173(clk,rst,matrix_A[6173],matrix_B[173],mul_res1[6173]);
multi_7x28 multi_7x28_mod_6174(clk,rst,matrix_A[6174],matrix_B[174],mul_res1[6174]);
multi_7x28 multi_7x28_mod_6175(clk,rst,matrix_A[6175],matrix_B[175],mul_res1[6175]);
multi_7x28 multi_7x28_mod_6176(clk,rst,matrix_A[6176],matrix_B[176],mul_res1[6176]);
multi_7x28 multi_7x28_mod_6177(clk,rst,matrix_A[6177],matrix_B[177],mul_res1[6177]);
multi_7x28 multi_7x28_mod_6178(clk,rst,matrix_A[6178],matrix_B[178],mul_res1[6178]);
multi_7x28 multi_7x28_mod_6179(clk,rst,matrix_A[6179],matrix_B[179],mul_res1[6179]);
multi_7x28 multi_7x28_mod_6180(clk,rst,matrix_A[6180],matrix_B[180],mul_res1[6180]);
multi_7x28 multi_7x28_mod_6181(clk,rst,matrix_A[6181],matrix_B[181],mul_res1[6181]);
multi_7x28 multi_7x28_mod_6182(clk,rst,matrix_A[6182],matrix_B[182],mul_res1[6182]);
multi_7x28 multi_7x28_mod_6183(clk,rst,matrix_A[6183],matrix_B[183],mul_res1[6183]);
multi_7x28 multi_7x28_mod_6184(clk,rst,matrix_A[6184],matrix_B[184],mul_res1[6184]);
multi_7x28 multi_7x28_mod_6185(clk,rst,matrix_A[6185],matrix_B[185],mul_res1[6185]);
multi_7x28 multi_7x28_mod_6186(clk,rst,matrix_A[6186],matrix_B[186],mul_res1[6186]);
multi_7x28 multi_7x28_mod_6187(clk,rst,matrix_A[6187],matrix_B[187],mul_res1[6187]);
multi_7x28 multi_7x28_mod_6188(clk,rst,matrix_A[6188],matrix_B[188],mul_res1[6188]);
multi_7x28 multi_7x28_mod_6189(clk,rst,matrix_A[6189],matrix_B[189],mul_res1[6189]);
multi_7x28 multi_7x28_mod_6190(clk,rst,matrix_A[6190],matrix_B[190],mul_res1[6190]);
multi_7x28 multi_7x28_mod_6191(clk,rst,matrix_A[6191],matrix_B[191],mul_res1[6191]);
multi_7x28 multi_7x28_mod_6192(clk,rst,matrix_A[6192],matrix_B[192],mul_res1[6192]);
multi_7x28 multi_7x28_mod_6193(clk,rst,matrix_A[6193],matrix_B[193],mul_res1[6193]);
multi_7x28 multi_7x28_mod_6194(clk,rst,matrix_A[6194],matrix_B[194],mul_res1[6194]);
multi_7x28 multi_7x28_mod_6195(clk,rst,matrix_A[6195],matrix_B[195],mul_res1[6195]);
multi_7x28 multi_7x28_mod_6196(clk,rst,matrix_A[6196],matrix_B[196],mul_res1[6196]);
multi_7x28 multi_7x28_mod_6197(clk,rst,matrix_A[6197],matrix_B[197],mul_res1[6197]);
multi_7x28 multi_7x28_mod_6198(clk,rst,matrix_A[6198],matrix_B[198],mul_res1[6198]);
multi_7x28 multi_7x28_mod_6199(clk,rst,matrix_A[6199],matrix_B[199],mul_res1[6199]);
multi_7x28 multi_7x28_mod_6200(clk,rst,matrix_A[6200],matrix_B[0],mul_res1[6200]);
multi_7x28 multi_7x28_mod_6201(clk,rst,matrix_A[6201],matrix_B[1],mul_res1[6201]);
multi_7x28 multi_7x28_mod_6202(clk,rst,matrix_A[6202],matrix_B[2],mul_res1[6202]);
multi_7x28 multi_7x28_mod_6203(clk,rst,matrix_A[6203],matrix_B[3],mul_res1[6203]);
multi_7x28 multi_7x28_mod_6204(clk,rst,matrix_A[6204],matrix_B[4],mul_res1[6204]);
multi_7x28 multi_7x28_mod_6205(clk,rst,matrix_A[6205],matrix_B[5],mul_res1[6205]);
multi_7x28 multi_7x28_mod_6206(clk,rst,matrix_A[6206],matrix_B[6],mul_res1[6206]);
multi_7x28 multi_7x28_mod_6207(clk,rst,matrix_A[6207],matrix_B[7],mul_res1[6207]);
multi_7x28 multi_7x28_mod_6208(clk,rst,matrix_A[6208],matrix_B[8],mul_res1[6208]);
multi_7x28 multi_7x28_mod_6209(clk,rst,matrix_A[6209],matrix_B[9],mul_res1[6209]);
multi_7x28 multi_7x28_mod_6210(clk,rst,matrix_A[6210],matrix_B[10],mul_res1[6210]);
multi_7x28 multi_7x28_mod_6211(clk,rst,matrix_A[6211],matrix_B[11],mul_res1[6211]);
multi_7x28 multi_7x28_mod_6212(clk,rst,matrix_A[6212],matrix_B[12],mul_res1[6212]);
multi_7x28 multi_7x28_mod_6213(clk,rst,matrix_A[6213],matrix_B[13],mul_res1[6213]);
multi_7x28 multi_7x28_mod_6214(clk,rst,matrix_A[6214],matrix_B[14],mul_res1[6214]);
multi_7x28 multi_7x28_mod_6215(clk,rst,matrix_A[6215],matrix_B[15],mul_res1[6215]);
multi_7x28 multi_7x28_mod_6216(clk,rst,matrix_A[6216],matrix_B[16],mul_res1[6216]);
multi_7x28 multi_7x28_mod_6217(clk,rst,matrix_A[6217],matrix_B[17],mul_res1[6217]);
multi_7x28 multi_7x28_mod_6218(clk,rst,matrix_A[6218],matrix_B[18],mul_res1[6218]);
multi_7x28 multi_7x28_mod_6219(clk,rst,matrix_A[6219],matrix_B[19],mul_res1[6219]);
multi_7x28 multi_7x28_mod_6220(clk,rst,matrix_A[6220],matrix_B[20],mul_res1[6220]);
multi_7x28 multi_7x28_mod_6221(clk,rst,matrix_A[6221],matrix_B[21],mul_res1[6221]);
multi_7x28 multi_7x28_mod_6222(clk,rst,matrix_A[6222],matrix_B[22],mul_res1[6222]);
multi_7x28 multi_7x28_mod_6223(clk,rst,matrix_A[6223],matrix_B[23],mul_res1[6223]);
multi_7x28 multi_7x28_mod_6224(clk,rst,matrix_A[6224],matrix_B[24],mul_res1[6224]);
multi_7x28 multi_7x28_mod_6225(clk,rst,matrix_A[6225],matrix_B[25],mul_res1[6225]);
multi_7x28 multi_7x28_mod_6226(clk,rst,matrix_A[6226],matrix_B[26],mul_res1[6226]);
multi_7x28 multi_7x28_mod_6227(clk,rst,matrix_A[6227],matrix_B[27],mul_res1[6227]);
multi_7x28 multi_7x28_mod_6228(clk,rst,matrix_A[6228],matrix_B[28],mul_res1[6228]);
multi_7x28 multi_7x28_mod_6229(clk,rst,matrix_A[6229],matrix_B[29],mul_res1[6229]);
multi_7x28 multi_7x28_mod_6230(clk,rst,matrix_A[6230],matrix_B[30],mul_res1[6230]);
multi_7x28 multi_7x28_mod_6231(clk,rst,matrix_A[6231],matrix_B[31],mul_res1[6231]);
multi_7x28 multi_7x28_mod_6232(clk,rst,matrix_A[6232],matrix_B[32],mul_res1[6232]);
multi_7x28 multi_7x28_mod_6233(clk,rst,matrix_A[6233],matrix_B[33],mul_res1[6233]);
multi_7x28 multi_7x28_mod_6234(clk,rst,matrix_A[6234],matrix_B[34],mul_res1[6234]);
multi_7x28 multi_7x28_mod_6235(clk,rst,matrix_A[6235],matrix_B[35],mul_res1[6235]);
multi_7x28 multi_7x28_mod_6236(clk,rst,matrix_A[6236],matrix_B[36],mul_res1[6236]);
multi_7x28 multi_7x28_mod_6237(clk,rst,matrix_A[6237],matrix_B[37],mul_res1[6237]);
multi_7x28 multi_7x28_mod_6238(clk,rst,matrix_A[6238],matrix_B[38],mul_res1[6238]);
multi_7x28 multi_7x28_mod_6239(clk,rst,matrix_A[6239],matrix_B[39],mul_res1[6239]);
multi_7x28 multi_7x28_mod_6240(clk,rst,matrix_A[6240],matrix_B[40],mul_res1[6240]);
multi_7x28 multi_7x28_mod_6241(clk,rst,matrix_A[6241],matrix_B[41],mul_res1[6241]);
multi_7x28 multi_7x28_mod_6242(clk,rst,matrix_A[6242],matrix_B[42],mul_res1[6242]);
multi_7x28 multi_7x28_mod_6243(clk,rst,matrix_A[6243],matrix_B[43],mul_res1[6243]);
multi_7x28 multi_7x28_mod_6244(clk,rst,matrix_A[6244],matrix_B[44],mul_res1[6244]);
multi_7x28 multi_7x28_mod_6245(clk,rst,matrix_A[6245],matrix_B[45],mul_res1[6245]);
multi_7x28 multi_7x28_mod_6246(clk,rst,matrix_A[6246],matrix_B[46],mul_res1[6246]);
multi_7x28 multi_7x28_mod_6247(clk,rst,matrix_A[6247],matrix_B[47],mul_res1[6247]);
multi_7x28 multi_7x28_mod_6248(clk,rst,matrix_A[6248],matrix_B[48],mul_res1[6248]);
multi_7x28 multi_7x28_mod_6249(clk,rst,matrix_A[6249],matrix_B[49],mul_res1[6249]);
multi_7x28 multi_7x28_mod_6250(clk,rst,matrix_A[6250],matrix_B[50],mul_res1[6250]);
multi_7x28 multi_7x28_mod_6251(clk,rst,matrix_A[6251],matrix_B[51],mul_res1[6251]);
multi_7x28 multi_7x28_mod_6252(clk,rst,matrix_A[6252],matrix_B[52],mul_res1[6252]);
multi_7x28 multi_7x28_mod_6253(clk,rst,matrix_A[6253],matrix_B[53],mul_res1[6253]);
multi_7x28 multi_7x28_mod_6254(clk,rst,matrix_A[6254],matrix_B[54],mul_res1[6254]);
multi_7x28 multi_7x28_mod_6255(clk,rst,matrix_A[6255],matrix_B[55],mul_res1[6255]);
multi_7x28 multi_7x28_mod_6256(clk,rst,matrix_A[6256],matrix_B[56],mul_res1[6256]);
multi_7x28 multi_7x28_mod_6257(clk,rst,matrix_A[6257],matrix_B[57],mul_res1[6257]);
multi_7x28 multi_7x28_mod_6258(clk,rst,matrix_A[6258],matrix_B[58],mul_res1[6258]);
multi_7x28 multi_7x28_mod_6259(clk,rst,matrix_A[6259],matrix_B[59],mul_res1[6259]);
multi_7x28 multi_7x28_mod_6260(clk,rst,matrix_A[6260],matrix_B[60],mul_res1[6260]);
multi_7x28 multi_7x28_mod_6261(clk,rst,matrix_A[6261],matrix_B[61],mul_res1[6261]);
multi_7x28 multi_7x28_mod_6262(clk,rst,matrix_A[6262],matrix_B[62],mul_res1[6262]);
multi_7x28 multi_7x28_mod_6263(clk,rst,matrix_A[6263],matrix_B[63],mul_res1[6263]);
multi_7x28 multi_7x28_mod_6264(clk,rst,matrix_A[6264],matrix_B[64],mul_res1[6264]);
multi_7x28 multi_7x28_mod_6265(clk,rst,matrix_A[6265],matrix_B[65],mul_res1[6265]);
multi_7x28 multi_7x28_mod_6266(clk,rst,matrix_A[6266],matrix_B[66],mul_res1[6266]);
multi_7x28 multi_7x28_mod_6267(clk,rst,matrix_A[6267],matrix_B[67],mul_res1[6267]);
multi_7x28 multi_7x28_mod_6268(clk,rst,matrix_A[6268],matrix_B[68],mul_res1[6268]);
multi_7x28 multi_7x28_mod_6269(clk,rst,matrix_A[6269],matrix_B[69],mul_res1[6269]);
multi_7x28 multi_7x28_mod_6270(clk,rst,matrix_A[6270],matrix_B[70],mul_res1[6270]);
multi_7x28 multi_7x28_mod_6271(clk,rst,matrix_A[6271],matrix_B[71],mul_res1[6271]);
multi_7x28 multi_7x28_mod_6272(clk,rst,matrix_A[6272],matrix_B[72],mul_res1[6272]);
multi_7x28 multi_7x28_mod_6273(clk,rst,matrix_A[6273],matrix_B[73],mul_res1[6273]);
multi_7x28 multi_7x28_mod_6274(clk,rst,matrix_A[6274],matrix_B[74],mul_res1[6274]);
multi_7x28 multi_7x28_mod_6275(clk,rst,matrix_A[6275],matrix_B[75],mul_res1[6275]);
multi_7x28 multi_7x28_mod_6276(clk,rst,matrix_A[6276],matrix_B[76],mul_res1[6276]);
multi_7x28 multi_7x28_mod_6277(clk,rst,matrix_A[6277],matrix_B[77],mul_res1[6277]);
multi_7x28 multi_7x28_mod_6278(clk,rst,matrix_A[6278],matrix_B[78],mul_res1[6278]);
multi_7x28 multi_7x28_mod_6279(clk,rst,matrix_A[6279],matrix_B[79],mul_res1[6279]);
multi_7x28 multi_7x28_mod_6280(clk,rst,matrix_A[6280],matrix_B[80],mul_res1[6280]);
multi_7x28 multi_7x28_mod_6281(clk,rst,matrix_A[6281],matrix_B[81],mul_res1[6281]);
multi_7x28 multi_7x28_mod_6282(clk,rst,matrix_A[6282],matrix_B[82],mul_res1[6282]);
multi_7x28 multi_7x28_mod_6283(clk,rst,matrix_A[6283],matrix_B[83],mul_res1[6283]);
multi_7x28 multi_7x28_mod_6284(clk,rst,matrix_A[6284],matrix_B[84],mul_res1[6284]);
multi_7x28 multi_7x28_mod_6285(clk,rst,matrix_A[6285],matrix_B[85],mul_res1[6285]);
multi_7x28 multi_7x28_mod_6286(clk,rst,matrix_A[6286],matrix_B[86],mul_res1[6286]);
multi_7x28 multi_7x28_mod_6287(clk,rst,matrix_A[6287],matrix_B[87],mul_res1[6287]);
multi_7x28 multi_7x28_mod_6288(clk,rst,matrix_A[6288],matrix_B[88],mul_res1[6288]);
multi_7x28 multi_7x28_mod_6289(clk,rst,matrix_A[6289],matrix_B[89],mul_res1[6289]);
multi_7x28 multi_7x28_mod_6290(clk,rst,matrix_A[6290],matrix_B[90],mul_res1[6290]);
multi_7x28 multi_7x28_mod_6291(clk,rst,matrix_A[6291],matrix_B[91],mul_res1[6291]);
multi_7x28 multi_7x28_mod_6292(clk,rst,matrix_A[6292],matrix_B[92],mul_res1[6292]);
multi_7x28 multi_7x28_mod_6293(clk,rst,matrix_A[6293],matrix_B[93],mul_res1[6293]);
multi_7x28 multi_7x28_mod_6294(clk,rst,matrix_A[6294],matrix_B[94],mul_res1[6294]);
multi_7x28 multi_7x28_mod_6295(clk,rst,matrix_A[6295],matrix_B[95],mul_res1[6295]);
multi_7x28 multi_7x28_mod_6296(clk,rst,matrix_A[6296],matrix_B[96],mul_res1[6296]);
multi_7x28 multi_7x28_mod_6297(clk,rst,matrix_A[6297],matrix_B[97],mul_res1[6297]);
multi_7x28 multi_7x28_mod_6298(clk,rst,matrix_A[6298],matrix_B[98],mul_res1[6298]);
multi_7x28 multi_7x28_mod_6299(clk,rst,matrix_A[6299],matrix_B[99],mul_res1[6299]);
multi_7x28 multi_7x28_mod_6300(clk,rst,matrix_A[6300],matrix_B[100],mul_res1[6300]);
multi_7x28 multi_7x28_mod_6301(clk,rst,matrix_A[6301],matrix_B[101],mul_res1[6301]);
multi_7x28 multi_7x28_mod_6302(clk,rst,matrix_A[6302],matrix_B[102],mul_res1[6302]);
multi_7x28 multi_7x28_mod_6303(clk,rst,matrix_A[6303],matrix_B[103],mul_res1[6303]);
multi_7x28 multi_7x28_mod_6304(clk,rst,matrix_A[6304],matrix_B[104],mul_res1[6304]);
multi_7x28 multi_7x28_mod_6305(clk,rst,matrix_A[6305],matrix_B[105],mul_res1[6305]);
multi_7x28 multi_7x28_mod_6306(clk,rst,matrix_A[6306],matrix_B[106],mul_res1[6306]);
multi_7x28 multi_7x28_mod_6307(clk,rst,matrix_A[6307],matrix_B[107],mul_res1[6307]);
multi_7x28 multi_7x28_mod_6308(clk,rst,matrix_A[6308],matrix_B[108],mul_res1[6308]);
multi_7x28 multi_7x28_mod_6309(clk,rst,matrix_A[6309],matrix_B[109],mul_res1[6309]);
multi_7x28 multi_7x28_mod_6310(clk,rst,matrix_A[6310],matrix_B[110],mul_res1[6310]);
multi_7x28 multi_7x28_mod_6311(clk,rst,matrix_A[6311],matrix_B[111],mul_res1[6311]);
multi_7x28 multi_7x28_mod_6312(clk,rst,matrix_A[6312],matrix_B[112],mul_res1[6312]);
multi_7x28 multi_7x28_mod_6313(clk,rst,matrix_A[6313],matrix_B[113],mul_res1[6313]);
multi_7x28 multi_7x28_mod_6314(clk,rst,matrix_A[6314],matrix_B[114],mul_res1[6314]);
multi_7x28 multi_7x28_mod_6315(clk,rst,matrix_A[6315],matrix_B[115],mul_res1[6315]);
multi_7x28 multi_7x28_mod_6316(clk,rst,matrix_A[6316],matrix_B[116],mul_res1[6316]);
multi_7x28 multi_7x28_mod_6317(clk,rst,matrix_A[6317],matrix_B[117],mul_res1[6317]);
multi_7x28 multi_7x28_mod_6318(clk,rst,matrix_A[6318],matrix_B[118],mul_res1[6318]);
multi_7x28 multi_7x28_mod_6319(clk,rst,matrix_A[6319],matrix_B[119],mul_res1[6319]);
multi_7x28 multi_7x28_mod_6320(clk,rst,matrix_A[6320],matrix_B[120],mul_res1[6320]);
multi_7x28 multi_7x28_mod_6321(clk,rst,matrix_A[6321],matrix_B[121],mul_res1[6321]);
multi_7x28 multi_7x28_mod_6322(clk,rst,matrix_A[6322],matrix_B[122],mul_res1[6322]);
multi_7x28 multi_7x28_mod_6323(clk,rst,matrix_A[6323],matrix_B[123],mul_res1[6323]);
multi_7x28 multi_7x28_mod_6324(clk,rst,matrix_A[6324],matrix_B[124],mul_res1[6324]);
multi_7x28 multi_7x28_mod_6325(clk,rst,matrix_A[6325],matrix_B[125],mul_res1[6325]);
multi_7x28 multi_7x28_mod_6326(clk,rst,matrix_A[6326],matrix_B[126],mul_res1[6326]);
multi_7x28 multi_7x28_mod_6327(clk,rst,matrix_A[6327],matrix_B[127],mul_res1[6327]);
multi_7x28 multi_7x28_mod_6328(clk,rst,matrix_A[6328],matrix_B[128],mul_res1[6328]);
multi_7x28 multi_7x28_mod_6329(clk,rst,matrix_A[6329],matrix_B[129],mul_res1[6329]);
multi_7x28 multi_7x28_mod_6330(clk,rst,matrix_A[6330],matrix_B[130],mul_res1[6330]);
multi_7x28 multi_7x28_mod_6331(clk,rst,matrix_A[6331],matrix_B[131],mul_res1[6331]);
multi_7x28 multi_7x28_mod_6332(clk,rst,matrix_A[6332],matrix_B[132],mul_res1[6332]);
multi_7x28 multi_7x28_mod_6333(clk,rst,matrix_A[6333],matrix_B[133],mul_res1[6333]);
multi_7x28 multi_7x28_mod_6334(clk,rst,matrix_A[6334],matrix_B[134],mul_res1[6334]);
multi_7x28 multi_7x28_mod_6335(clk,rst,matrix_A[6335],matrix_B[135],mul_res1[6335]);
multi_7x28 multi_7x28_mod_6336(clk,rst,matrix_A[6336],matrix_B[136],mul_res1[6336]);
multi_7x28 multi_7x28_mod_6337(clk,rst,matrix_A[6337],matrix_B[137],mul_res1[6337]);
multi_7x28 multi_7x28_mod_6338(clk,rst,matrix_A[6338],matrix_B[138],mul_res1[6338]);
multi_7x28 multi_7x28_mod_6339(clk,rst,matrix_A[6339],matrix_B[139],mul_res1[6339]);
multi_7x28 multi_7x28_mod_6340(clk,rst,matrix_A[6340],matrix_B[140],mul_res1[6340]);
multi_7x28 multi_7x28_mod_6341(clk,rst,matrix_A[6341],matrix_B[141],mul_res1[6341]);
multi_7x28 multi_7x28_mod_6342(clk,rst,matrix_A[6342],matrix_B[142],mul_res1[6342]);
multi_7x28 multi_7x28_mod_6343(clk,rst,matrix_A[6343],matrix_B[143],mul_res1[6343]);
multi_7x28 multi_7x28_mod_6344(clk,rst,matrix_A[6344],matrix_B[144],mul_res1[6344]);
multi_7x28 multi_7x28_mod_6345(clk,rst,matrix_A[6345],matrix_B[145],mul_res1[6345]);
multi_7x28 multi_7x28_mod_6346(clk,rst,matrix_A[6346],matrix_B[146],mul_res1[6346]);
multi_7x28 multi_7x28_mod_6347(clk,rst,matrix_A[6347],matrix_B[147],mul_res1[6347]);
multi_7x28 multi_7x28_mod_6348(clk,rst,matrix_A[6348],matrix_B[148],mul_res1[6348]);
multi_7x28 multi_7x28_mod_6349(clk,rst,matrix_A[6349],matrix_B[149],mul_res1[6349]);
multi_7x28 multi_7x28_mod_6350(clk,rst,matrix_A[6350],matrix_B[150],mul_res1[6350]);
multi_7x28 multi_7x28_mod_6351(clk,rst,matrix_A[6351],matrix_B[151],mul_res1[6351]);
multi_7x28 multi_7x28_mod_6352(clk,rst,matrix_A[6352],matrix_B[152],mul_res1[6352]);
multi_7x28 multi_7x28_mod_6353(clk,rst,matrix_A[6353],matrix_B[153],mul_res1[6353]);
multi_7x28 multi_7x28_mod_6354(clk,rst,matrix_A[6354],matrix_B[154],mul_res1[6354]);
multi_7x28 multi_7x28_mod_6355(clk,rst,matrix_A[6355],matrix_B[155],mul_res1[6355]);
multi_7x28 multi_7x28_mod_6356(clk,rst,matrix_A[6356],matrix_B[156],mul_res1[6356]);
multi_7x28 multi_7x28_mod_6357(clk,rst,matrix_A[6357],matrix_B[157],mul_res1[6357]);
multi_7x28 multi_7x28_mod_6358(clk,rst,matrix_A[6358],matrix_B[158],mul_res1[6358]);
multi_7x28 multi_7x28_mod_6359(clk,rst,matrix_A[6359],matrix_B[159],mul_res1[6359]);
multi_7x28 multi_7x28_mod_6360(clk,rst,matrix_A[6360],matrix_B[160],mul_res1[6360]);
multi_7x28 multi_7x28_mod_6361(clk,rst,matrix_A[6361],matrix_B[161],mul_res1[6361]);
multi_7x28 multi_7x28_mod_6362(clk,rst,matrix_A[6362],matrix_B[162],mul_res1[6362]);
multi_7x28 multi_7x28_mod_6363(clk,rst,matrix_A[6363],matrix_B[163],mul_res1[6363]);
multi_7x28 multi_7x28_mod_6364(clk,rst,matrix_A[6364],matrix_B[164],mul_res1[6364]);
multi_7x28 multi_7x28_mod_6365(clk,rst,matrix_A[6365],matrix_B[165],mul_res1[6365]);
multi_7x28 multi_7x28_mod_6366(clk,rst,matrix_A[6366],matrix_B[166],mul_res1[6366]);
multi_7x28 multi_7x28_mod_6367(clk,rst,matrix_A[6367],matrix_B[167],mul_res1[6367]);
multi_7x28 multi_7x28_mod_6368(clk,rst,matrix_A[6368],matrix_B[168],mul_res1[6368]);
multi_7x28 multi_7x28_mod_6369(clk,rst,matrix_A[6369],matrix_B[169],mul_res1[6369]);
multi_7x28 multi_7x28_mod_6370(clk,rst,matrix_A[6370],matrix_B[170],mul_res1[6370]);
multi_7x28 multi_7x28_mod_6371(clk,rst,matrix_A[6371],matrix_B[171],mul_res1[6371]);
multi_7x28 multi_7x28_mod_6372(clk,rst,matrix_A[6372],matrix_B[172],mul_res1[6372]);
multi_7x28 multi_7x28_mod_6373(clk,rst,matrix_A[6373],matrix_B[173],mul_res1[6373]);
multi_7x28 multi_7x28_mod_6374(clk,rst,matrix_A[6374],matrix_B[174],mul_res1[6374]);
multi_7x28 multi_7x28_mod_6375(clk,rst,matrix_A[6375],matrix_B[175],mul_res1[6375]);
multi_7x28 multi_7x28_mod_6376(clk,rst,matrix_A[6376],matrix_B[176],mul_res1[6376]);
multi_7x28 multi_7x28_mod_6377(clk,rst,matrix_A[6377],matrix_B[177],mul_res1[6377]);
multi_7x28 multi_7x28_mod_6378(clk,rst,matrix_A[6378],matrix_B[178],mul_res1[6378]);
multi_7x28 multi_7x28_mod_6379(clk,rst,matrix_A[6379],matrix_B[179],mul_res1[6379]);
multi_7x28 multi_7x28_mod_6380(clk,rst,matrix_A[6380],matrix_B[180],mul_res1[6380]);
multi_7x28 multi_7x28_mod_6381(clk,rst,matrix_A[6381],matrix_B[181],mul_res1[6381]);
multi_7x28 multi_7x28_mod_6382(clk,rst,matrix_A[6382],matrix_B[182],mul_res1[6382]);
multi_7x28 multi_7x28_mod_6383(clk,rst,matrix_A[6383],matrix_B[183],mul_res1[6383]);
multi_7x28 multi_7x28_mod_6384(clk,rst,matrix_A[6384],matrix_B[184],mul_res1[6384]);
multi_7x28 multi_7x28_mod_6385(clk,rst,matrix_A[6385],matrix_B[185],mul_res1[6385]);
multi_7x28 multi_7x28_mod_6386(clk,rst,matrix_A[6386],matrix_B[186],mul_res1[6386]);
multi_7x28 multi_7x28_mod_6387(clk,rst,matrix_A[6387],matrix_B[187],mul_res1[6387]);
multi_7x28 multi_7x28_mod_6388(clk,rst,matrix_A[6388],matrix_B[188],mul_res1[6388]);
multi_7x28 multi_7x28_mod_6389(clk,rst,matrix_A[6389],matrix_B[189],mul_res1[6389]);
multi_7x28 multi_7x28_mod_6390(clk,rst,matrix_A[6390],matrix_B[190],mul_res1[6390]);
multi_7x28 multi_7x28_mod_6391(clk,rst,matrix_A[6391],matrix_B[191],mul_res1[6391]);
multi_7x28 multi_7x28_mod_6392(clk,rst,matrix_A[6392],matrix_B[192],mul_res1[6392]);
multi_7x28 multi_7x28_mod_6393(clk,rst,matrix_A[6393],matrix_B[193],mul_res1[6393]);
multi_7x28 multi_7x28_mod_6394(clk,rst,matrix_A[6394],matrix_B[194],mul_res1[6394]);
multi_7x28 multi_7x28_mod_6395(clk,rst,matrix_A[6395],matrix_B[195],mul_res1[6395]);
multi_7x28 multi_7x28_mod_6396(clk,rst,matrix_A[6396],matrix_B[196],mul_res1[6396]);
multi_7x28 multi_7x28_mod_6397(clk,rst,matrix_A[6397],matrix_B[197],mul_res1[6397]);
multi_7x28 multi_7x28_mod_6398(clk,rst,matrix_A[6398],matrix_B[198],mul_res1[6398]);
multi_7x28 multi_7x28_mod_6399(clk,rst,matrix_A[6399],matrix_B[199],mul_res1[6399]);
multi_7x28 multi_7x28_mod_6400(clk,rst,matrix_A[6400],matrix_B[0],mul_res1[6400]);
multi_7x28 multi_7x28_mod_6401(clk,rst,matrix_A[6401],matrix_B[1],mul_res1[6401]);
multi_7x28 multi_7x28_mod_6402(clk,rst,matrix_A[6402],matrix_B[2],mul_res1[6402]);
multi_7x28 multi_7x28_mod_6403(clk,rst,matrix_A[6403],matrix_B[3],mul_res1[6403]);
multi_7x28 multi_7x28_mod_6404(clk,rst,matrix_A[6404],matrix_B[4],mul_res1[6404]);
multi_7x28 multi_7x28_mod_6405(clk,rst,matrix_A[6405],matrix_B[5],mul_res1[6405]);
multi_7x28 multi_7x28_mod_6406(clk,rst,matrix_A[6406],matrix_B[6],mul_res1[6406]);
multi_7x28 multi_7x28_mod_6407(clk,rst,matrix_A[6407],matrix_B[7],mul_res1[6407]);
multi_7x28 multi_7x28_mod_6408(clk,rst,matrix_A[6408],matrix_B[8],mul_res1[6408]);
multi_7x28 multi_7x28_mod_6409(clk,rst,matrix_A[6409],matrix_B[9],mul_res1[6409]);
multi_7x28 multi_7x28_mod_6410(clk,rst,matrix_A[6410],matrix_B[10],mul_res1[6410]);
multi_7x28 multi_7x28_mod_6411(clk,rst,matrix_A[6411],matrix_B[11],mul_res1[6411]);
multi_7x28 multi_7x28_mod_6412(clk,rst,matrix_A[6412],matrix_B[12],mul_res1[6412]);
multi_7x28 multi_7x28_mod_6413(clk,rst,matrix_A[6413],matrix_B[13],mul_res1[6413]);
multi_7x28 multi_7x28_mod_6414(clk,rst,matrix_A[6414],matrix_B[14],mul_res1[6414]);
multi_7x28 multi_7x28_mod_6415(clk,rst,matrix_A[6415],matrix_B[15],mul_res1[6415]);
multi_7x28 multi_7x28_mod_6416(clk,rst,matrix_A[6416],matrix_B[16],mul_res1[6416]);
multi_7x28 multi_7x28_mod_6417(clk,rst,matrix_A[6417],matrix_B[17],mul_res1[6417]);
multi_7x28 multi_7x28_mod_6418(clk,rst,matrix_A[6418],matrix_B[18],mul_res1[6418]);
multi_7x28 multi_7x28_mod_6419(clk,rst,matrix_A[6419],matrix_B[19],mul_res1[6419]);
multi_7x28 multi_7x28_mod_6420(clk,rst,matrix_A[6420],matrix_B[20],mul_res1[6420]);
multi_7x28 multi_7x28_mod_6421(clk,rst,matrix_A[6421],matrix_B[21],mul_res1[6421]);
multi_7x28 multi_7x28_mod_6422(clk,rst,matrix_A[6422],matrix_B[22],mul_res1[6422]);
multi_7x28 multi_7x28_mod_6423(clk,rst,matrix_A[6423],matrix_B[23],mul_res1[6423]);
multi_7x28 multi_7x28_mod_6424(clk,rst,matrix_A[6424],matrix_B[24],mul_res1[6424]);
multi_7x28 multi_7x28_mod_6425(clk,rst,matrix_A[6425],matrix_B[25],mul_res1[6425]);
multi_7x28 multi_7x28_mod_6426(clk,rst,matrix_A[6426],matrix_B[26],mul_res1[6426]);
multi_7x28 multi_7x28_mod_6427(clk,rst,matrix_A[6427],matrix_B[27],mul_res1[6427]);
multi_7x28 multi_7x28_mod_6428(clk,rst,matrix_A[6428],matrix_B[28],mul_res1[6428]);
multi_7x28 multi_7x28_mod_6429(clk,rst,matrix_A[6429],matrix_B[29],mul_res1[6429]);
multi_7x28 multi_7x28_mod_6430(clk,rst,matrix_A[6430],matrix_B[30],mul_res1[6430]);
multi_7x28 multi_7x28_mod_6431(clk,rst,matrix_A[6431],matrix_B[31],mul_res1[6431]);
multi_7x28 multi_7x28_mod_6432(clk,rst,matrix_A[6432],matrix_B[32],mul_res1[6432]);
multi_7x28 multi_7x28_mod_6433(clk,rst,matrix_A[6433],matrix_B[33],mul_res1[6433]);
multi_7x28 multi_7x28_mod_6434(clk,rst,matrix_A[6434],matrix_B[34],mul_res1[6434]);
multi_7x28 multi_7x28_mod_6435(clk,rst,matrix_A[6435],matrix_B[35],mul_res1[6435]);
multi_7x28 multi_7x28_mod_6436(clk,rst,matrix_A[6436],matrix_B[36],mul_res1[6436]);
multi_7x28 multi_7x28_mod_6437(clk,rst,matrix_A[6437],matrix_B[37],mul_res1[6437]);
multi_7x28 multi_7x28_mod_6438(clk,rst,matrix_A[6438],matrix_B[38],mul_res1[6438]);
multi_7x28 multi_7x28_mod_6439(clk,rst,matrix_A[6439],matrix_B[39],mul_res1[6439]);
multi_7x28 multi_7x28_mod_6440(clk,rst,matrix_A[6440],matrix_B[40],mul_res1[6440]);
multi_7x28 multi_7x28_mod_6441(clk,rst,matrix_A[6441],matrix_B[41],mul_res1[6441]);
multi_7x28 multi_7x28_mod_6442(clk,rst,matrix_A[6442],matrix_B[42],mul_res1[6442]);
multi_7x28 multi_7x28_mod_6443(clk,rst,matrix_A[6443],matrix_B[43],mul_res1[6443]);
multi_7x28 multi_7x28_mod_6444(clk,rst,matrix_A[6444],matrix_B[44],mul_res1[6444]);
multi_7x28 multi_7x28_mod_6445(clk,rst,matrix_A[6445],matrix_B[45],mul_res1[6445]);
multi_7x28 multi_7x28_mod_6446(clk,rst,matrix_A[6446],matrix_B[46],mul_res1[6446]);
multi_7x28 multi_7x28_mod_6447(clk,rst,matrix_A[6447],matrix_B[47],mul_res1[6447]);
multi_7x28 multi_7x28_mod_6448(clk,rst,matrix_A[6448],matrix_B[48],mul_res1[6448]);
multi_7x28 multi_7x28_mod_6449(clk,rst,matrix_A[6449],matrix_B[49],mul_res1[6449]);
multi_7x28 multi_7x28_mod_6450(clk,rst,matrix_A[6450],matrix_B[50],mul_res1[6450]);
multi_7x28 multi_7x28_mod_6451(clk,rst,matrix_A[6451],matrix_B[51],mul_res1[6451]);
multi_7x28 multi_7x28_mod_6452(clk,rst,matrix_A[6452],matrix_B[52],mul_res1[6452]);
multi_7x28 multi_7x28_mod_6453(clk,rst,matrix_A[6453],matrix_B[53],mul_res1[6453]);
multi_7x28 multi_7x28_mod_6454(clk,rst,matrix_A[6454],matrix_B[54],mul_res1[6454]);
multi_7x28 multi_7x28_mod_6455(clk,rst,matrix_A[6455],matrix_B[55],mul_res1[6455]);
multi_7x28 multi_7x28_mod_6456(clk,rst,matrix_A[6456],matrix_B[56],mul_res1[6456]);
multi_7x28 multi_7x28_mod_6457(clk,rst,matrix_A[6457],matrix_B[57],mul_res1[6457]);
multi_7x28 multi_7x28_mod_6458(clk,rst,matrix_A[6458],matrix_B[58],mul_res1[6458]);
multi_7x28 multi_7x28_mod_6459(clk,rst,matrix_A[6459],matrix_B[59],mul_res1[6459]);
multi_7x28 multi_7x28_mod_6460(clk,rst,matrix_A[6460],matrix_B[60],mul_res1[6460]);
multi_7x28 multi_7x28_mod_6461(clk,rst,matrix_A[6461],matrix_B[61],mul_res1[6461]);
multi_7x28 multi_7x28_mod_6462(clk,rst,matrix_A[6462],matrix_B[62],mul_res1[6462]);
multi_7x28 multi_7x28_mod_6463(clk,rst,matrix_A[6463],matrix_B[63],mul_res1[6463]);
multi_7x28 multi_7x28_mod_6464(clk,rst,matrix_A[6464],matrix_B[64],mul_res1[6464]);
multi_7x28 multi_7x28_mod_6465(clk,rst,matrix_A[6465],matrix_B[65],mul_res1[6465]);
multi_7x28 multi_7x28_mod_6466(clk,rst,matrix_A[6466],matrix_B[66],mul_res1[6466]);
multi_7x28 multi_7x28_mod_6467(clk,rst,matrix_A[6467],matrix_B[67],mul_res1[6467]);
multi_7x28 multi_7x28_mod_6468(clk,rst,matrix_A[6468],matrix_B[68],mul_res1[6468]);
multi_7x28 multi_7x28_mod_6469(clk,rst,matrix_A[6469],matrix_B[69],mul_res1[6469]);
multi_7x28 multi_7x28_mod_6470(clk,rst,matrix_A[6470],matrix_B[70],mul_res1[6470]);
multi_7x28 multi_7x28_mod_6471(clk,rst,matrix_A[6471],matrix_B[71],mul_res1[6471]);
multi_7x28 multi_7x28_mod_6472(clk,rst,matrix_A[6472],matrix_B[72],mul_res1[6472]);
multi_7x28 multi_7x28_mod_6473(clk,rst,matrix_A[6473],matrix_B[73],mul_res1[6473]);
multi_7x28 multi_7x28_mod_6474(clk,rst,matrix_A[6474],matrix_B[74],mul_res1[6474]);
multi_7x28 multi_7x28_mod_6475(clk,rst,matrix_A[6475],matrix_B[75],mul_res1[6475]);
multi_7x28 multi_7x28_mod_6476(clk,rst,matrix_A[6476],matrix_B[76],mul_res1[6476]);
multi_7x28 multi_7x28_mod_6477(clk,rst,matrix_A[6477],matrix_B[77],mul_res1[6477]);
multi_7x28 multi_7x28_mod_6478(clk,rst,matrix_A[6478],matrix_B[78],mul_res1[6478]);
multi_7x28 multi_7x28_mod_6479(clk,rst,matrix_A[6479],matrix_B[79],mul_res1[6479]);
multi_7x28 multi_7x28_mod_6480(clk,rst,matrix_A[6480],matrix_B[80],mul_res1[6480]);
multi_7x28 multi_7x28_mod_6481(clk,rst,matrix_A[6481],matrix_B[81],mul_res1[6481]);
multi_7x28 multi_7x28_mod_6482(clk,rst,matrix_A[6482],matrix_B[82],mul_res1[6482]);
multi_7x28 multi_7x28_mod_6483(clk,rst,matrix_A[6483],matrix_B[83],mul_res1[6483]);
multi_7x28 multi_7x28_mod_6484(clk,rst,matrix_A[6484],matrix_B[84],mul_res1[6484]);
multi_7x28 multi_7x28_mod_6485(clk,rst,matrix_A[6485],matrix_B[85],mul_res1[6485]);
multi_7x28 multi_7x28_mod_6486(clk,rst,matrix_A[6486],matrix_B[86],mul_res1[6486]);
multi_7x28 multi_7x28_mod_6487(clk,rst,matrix_A[6487],matrix_B[87],mul_res1[6487]);
multi_7x28 multi_7x28_mod_6488(clk,rst,matrix_A[6488],matrix_B[88],mul_res1[6488]);
multi_7x28 multi_7x28_mod_6489(clk,rst,matrix_A[6489],matrix_B[89],mul_res1[6489]);
multi_7x28 multi_7x28_mod_6490(clk,rst,matrix_A[6490],matrix_B[90],mul_res1[6490]);
multi_7x28 multi_7x28_mod_6491(clk,rst,matrix_A[6491],matrix_B[91],mul_res1[6491]);
multi_7x28 multi_7x28_mod_6492(clk,rst,matrix_A[6492],matrix_B[92],mul_res1[6492]);
multi_7x28 multi_7x28_mod_6493(clk,rst,matrix_A[6493],matrix_B[93],mul_res1[6493]);
multi_7x28 multi_7x28_mod_6494(clk,rst,matrix_A[6494],matrix_B[94],mul_res1[6494]);
multi_7x28 multi_7x28_mod_6495(clk,rst,matrix_A[6495],matrix_B[95],mul_res1[6495]);
multi_7x28 multi_7x28_mod_6496(clk,rst,matrix_A[6496],matrix_B[96],mul_res1[6496]);
multi_7x28 multi_7x28_mod_6497(clk,rst,matrix_A[6497],matrix_B[97],mul_res1[6497]);
multi_7x28 multi_7x28_mod_6498(clk,rst,matrix_A[6498],matrix_B[98],mul_res1[6498]);
multi_7x28 multi_7x28_mod_6499(clk,rst,matrix_A[6499],matrix_B[99],mul_res1[6499]);
multi_7x28 multi_7x28_mod_6500(clk,rst,matrix_A[6500],matrix_B[100],mul_res1[6500]);
multi_7x28 multi_7x28_mod_6501(clk,rst,matrix_A[6501],matrix_B[101],mul_res1[6501]);
multi_7x28 multi_7x28_mod_6502(clk,rst,matrix_A[6502],matrix_B[102],mul_res1[6502]);
multi_7x28 multi_7x28_mod_6503(clk,rst,matrix_A[6503],matrix_B[103],mul_res1[6503]);
multi_7x28 multi_7x28_mod_6504(clk,rst,matrix_A[6504],matrix_B[104],mul_res1[6504]);
multi_7x28 multi_7x28_mod_6505(clk,rst,matrix_A[6505],matrix_B[105],mul_res1[6505]);
multi_7x28 multi_7x28_mod_6506(clk,rst,matrix_A[6506],matrix_B[106],mul_res1[6506]);
multi_7x28 multi_7x28_mod_6507(clk,rst,matrix_A[6507],matrix_B[107],mul_res1[6507]);
multi_7x28 multi_7x28_mod_6508(clk,rst,matrix_A[6508],matrix_B[108],mul_res1[6508]);
multi_7x28 multi_7x28_mod_6509(clk,rst,matrix_A[6509],matrix_B[109],mul_res1[6509]);
multi_7x28 multi_7x28_mod_6510(clk,rst,matrix_A[6510],matrix_B[110],mul_res1[6510]);
multi_7x28 multi_7x28_mod_6511(clk,rst,matrix_A[6511],matrix_B[111],mul_res1[6511]);
multi_7x28 multi_7x28_mod_6512(clk,rst,matrix_A[6512],matrix_B[112],mul_res1[6512]);
multi_7x28 multi_7x28_mod_6513(clk,rst,matrix_A[6513],matrix_B[113],mul_res1[6513]);
multi_7x28 multi_7x28_mod_6514(clk,rst,matrix_A[6514],matrix_B[114],mul_res1[6514]);
multi_7x28 multi_7x28_mod_6515(clk,rst,matrix_A[6515],matrix_B[115],mul_res1[6515]);
multi_7x28 multi_7x28_mod_6516(clk,rst,matrix_A[6516],matrix_B[116],mul_res1[6516]);
multi_7x28 multi_7x28_mod_6517(clk,rst,matrix_A[6517],matrix_B[117],mul_res1[6517]);
multi_7x28 multi_7x28_mod_6518(clk,rst,matrix_A[6518],matrix_B[118],mul_res1[6518]);
multi_7x28 multi_7x28_mod_6519(clk,rst,matrix_A[6519],matrix_B[119],mul_res1[6519]);
multi_7x28 multi_7x28_mod_6520(clk,rst,matrix_A[6520],matrix_B[120],mul_res1[6520]);
multi_7x28 multi_7x28_mod_6521(clk,rst,matrix_A[6521],matrix_B[121],mul_res1[6521]);
multi_7x28 multi_7x28_mod_6522(clk,rst,matrix_A[6522],matrix_B[122],mul_res1[6522]);
multi_7x28 multi_7x28_mod_6523(clk,rst,matrix_A[6523],matrix_B[123],mul_res1[6523]);
multi_7x28 multi_7x28_mod_6524(clk,rst,matrix_A[6524],matrix_B[124],mul_res1[6524]);
multi_7x28 multi_7x28_mod_6525(clk,rst,matrix_A[6525],matrix_B[125],mul_res1[6525]);
multi_7x28 multi_7x28_mod_6526(clk,rst,matrix_A[6526],matrix_B[126],mul_res1[6526]);
multi_7x28 multi_7x28_mod_6527(clk,rst,matrix_A[6527],matrix_B[127],mul_res1[6527]);
multi_7x28 multi_7x28_mod_6528(clk,rst,matrix_A[6528],matrix_B[128],mul_res1[6528]);
multi_7x28 multi_7x28_mod_6529(clk,rst,matrix_A[6529],matrix_B[129],mul_res1[6529]);
multi_7x28 multi_7x28_mod_6530(clk,rst,matrix_A[6530],matrix_B[130],mul_res1[6530]);
multi_7x28 multi_7x28_mod_6531(clk,rst,matrix_A[6531],matrix_B[131],mul_res1[6531]);
multi_7x28 multi_7x28_mod_6532(clk,rst,matrix_A[6532],matrix_B[132],mul_res1[6532]);
multi_7x28 multi_7x28_mod_6533(clk,rst,matrix_A[6533],matrix_B[133],mul_res1[6533]);
multi_7x28 multi_7x28_mod_6534(clk,rst,matrix_A[6534],matrix_B[134],mul_res1[6534]);
multi_7x28 multi_7x28_mod_6535(clk,rst,matrix_A[6535],matrix_B[135],mul_res1[6535]);
multi_7x28 multi_7x28_mod_6536(clk,rst,matrix_A[6536],matrix_B[136],mul_res1[6536]);
multi_7x28 multi_7x28_mod_6537(clk,rst,matrix_A[6537],matrix_B[137],mul_res1[6537]);
multi_7x28 multi_7x28_mod_6538(clk,rst,matrix_A[6538],matrix_B[138],mul_res1[6538]);
multi_7x28 multi_7x28_mod_6539(clk,rst,matrix_A[6539],matrix_B[139],mul_res1[6539]);
multi_7x28 multi_7x28_mod_6540(clk,rst,matrix_A[6540],matrix_B[140],mul_res1[6540]);
multi_7x28 multi_7x28_mod_6541(clk,rst,matrix_A[6541],matrix_B[141],mul_res1[6541]);
multi_7x28 multi_7x28_mod_6542(clk,rst,matrix_A[6542],matrix_B[142],mul_res1[6542]);
multi_7x28 multi_7x28_mod_6543(clk,rst,matrix_A[6543],matrix_B[143],mul_res1[6543]);
multi_7x28 multi_7x28_mod_6544(clk,rst,matrix_A[6544],matrix_B[144],mul_res1[6544]);
multi_7x28 multi_7x28_mod_6545(clk,rst,matrix_A[6545],matrix_B[145],mul_res1[6545]);
multi_7x28 multi_7x28_mod_6546(clk,rst,matrix_A[6546],matrix_B[146],mul_res1[6546]);
multi_7x28 multi_7x28_mod_6547(clk,rst,matrix_A[6547],matrix_B[147],mul_res1[6547]);
multi_7x28 multi_7x28_mod_6548(clk,rst,matrix_A[6548],matrix_B[148],mul_res1[6548]);
multi_7x28 multi_7x28_mod_6549(clk,rst,matrix_A[6549],matrix_B[149],mul_res1[6549]);
multi_7x28 multi_7x28_mod_6550(clk,rst,matrix_A[6550],matrix_B[150],mul_res1[6550]);
multi_7x28 multi_7x28_mod_6551(clk,rst,matrix_A[6551],matrix_B[151],mul_res1[6551]);
multi_7x28 multi_7x28_mod_6552(clk,rst,matrix_A[6552],matrix_B[152],mul_res1[6552]);
multi_7x28 multi_7x28_mod_6553(clk,rst,matrix_A[6553],matrix_B[153],mul_res1[6553]);
multi_7x28 multi_7x28_mod_6554(clk,rst,matrix_A[6554],matrix_B[154],mul_res1[6554]);
multi_7x28 multi_7x28_mod_6555(clk,rst,matrix_A[6555],matrix_B[155],mul_res1[6555]);
multi_7x28 multi_7x28_mod_6556(clk,rst,matrix_A[6556],matrix_B[156],mul_res1[6556]);
multi_7x28 multi_7x28_mod_6557(clk,rst,matrix_A[6557],matrix_B[157],mul_res1[6557]);
multi_7x28 multi_7x28_mod_6558(clk,rst,matrix_A[6558],matrix_B[158],mul_res1[6558]);
multi_7x28 multi_7x28_mod_6559(clk,rst,matrix_A[6559],matrix_B[159],mul_res1[6559]);
multi_7x28 multi_7x28_mod_6560(clk,rst,matrix_A[6560],matrix_B[160],mul_res1[6560]);
multi_7x28 multi_7x28_mod_6561(clk,rst,matrix_A[6561],matrix_B[161],mul_res1[6561]);
multi_7x28 multi_7x28_mod_6562(clk,rst,matrix_A[6562],matrix_B[162],mul_res1[6562]);
multi_7x28 multi_7x28_mod_6563(clk,rst,matrix_A[6563],matrix_B[163],mul_res1[6563]);
multi_7x28 multi_7x28_mod_6564(clk,rst,matrix_A[6564],matrix_B[164],mul_res1[6564]);
multi_7x28 multi_7x28_mod_6565(clk,rst,matrix_A[6565],matrix_B[165],mul_res1[6565]);
multi_7x28 multi_7x28_mod_6566(clk,rst,matrix_A[6566],matrix_B[166],mul_res1[6566]);
multi_7x28 multi_7x28_mod_6567(clk,rst,matrix_A[6567],matrix_B[167],mul_res1[6567]);
multi_7x28 multi_7x28_mod_6568(clk,rst,matrix_A[6568],matrix_B[168],mul_res1[6568]);
multi_7x28 multi_7x28_mod_6569(clk,rst,matrix_A[6569],matrix_B[169],mul_res1[6569]);
multi_7x28 multi_7x28_mod_6570(clk,rst,matrix_A[6570],matrix_B[170],mul_res1[6570]);
multi_7x28 multi_7x28_mod_6571(clk,rst,matrix_A[6571],matrix_B[171],mul_res1[6571]);
multi_7x28 multi_7x28_mod_6572(clk,rst,matrix_A[6572],matrix_B[172],mul_res1[6572]);
multi_7x28 multi_7x28_mod_6573(clk,rst,matrix_A[6573],matrix_B[173],mul_res1[6573]);
multi_7x28 multi_7x28_mod_6574(clk,rst,matrix_A[6574],matrix_B[174],mul_res1[6574]);
multi_7x28 multi_7x28_mod_6575(clk,rst,matrix_A[6575],matrix_B[175],mul_res1[6575]);
multi_7x28 multi_7x28_mod_6576(clk,rst,matrix_A[6576],matrix_B[176],mul_res1[6576]);
multi_7x28 multi_7x28_mod_6577(clk,rst,matrix_A[6577],matrix_B[177],mul_res1[6577]);
multi_7x28 multi_7x28_mod_6578(clk,rst,matrix_A[6578],matrix_B[178],mul_res1[6578]);
multi_7x28 multi_7x28_mod_6579(clk,rst,matrix_A[6579],matrix_B[179],mul_res1[6579]);
multi_7x28 multi_7x28_mod_6580(clk,rst,matrix_A[6580],matrix_B[180],mul_res1[6580]);
multi_7x28 multi_7x28_mod_6581(clk,rst,matrix_A[6581],matrix_B[181],mul_res1[6581]);
multi_7x28 multi_7x28_mod_6582(clk,rst,matrix_A[6582],matrix_B[182],mul_res1[6582]);
multi_7x28 multi_7x28_mod_6583(clk,rst,matrix_A[6583],matrix_B[183],mul_res1[6583]);
multi_7x28 multi_7x28_mod_6584(clk,rst,matrix_A[6584],matrix_B[184],mul_res1[6584]);
multi_7x28 multi_7x28_mod_6585(clk,rst,matrix_A[6585],matrix_B[185],mul_res1[6585]);
multi_7x28 multi_7x28_mod_6586(clk,rst,matrix_A[6586],matrix_B[186],mul_res1[6586]);
multi_7x28 multi_7x28_mod_6587(clk,rst,matrix_A[6587],matrix_B[187],mul_res1[6587]);
multi_7x28 multi_7x28_mod_6588(clk,rst,matrix_A[6588],matrix_B[188],mul_res1[6588]);
multi_7x28 multi_7x28_mod_6589(clk,rst,matrix_A[6589],matrix_B[189],mul_res1[6589]);
multi_7x28 multi_7x28_mod_6590(clk,rst,matrix_A[6590],matrix_B[190],mul_res1[6590]);
multi_7x28 multi_7x28_mod_6591(clk,rst,matrix_A[6591],matrix_B[191],mul_res1[6591]);
multi_7x28 multi_7x28_mod_6592(clk,rst,matrix_A[6592],matrix_B[192],mul_res1[6592]);
multi_7x28 multi_7x28_mod_6593(clk,rst,matrix_A[6593],matrix_B[193],mul_res1[6593]);
multi_7x28 multi_7x28_mod_6594(clk,rst,matrix_A[6594],matrix_B[194],mul_res1[6594]);
multi_7x28 multi_7x28_mod_6595(clk,rst,matrix_A[6595],matrix_B[195],mul_res1[6595]);
multi_7x28 multi_7x28_mod_6596(clk,rst,matrix_A[6596],matrix_B[196],mul_res1[6596]);
multi_7x28 multi_7x28_mod_6597(clk,rst,matrix_A[6597],matrix_B[197],mul_res1[6597]);
multi_7x28 multi_7x28_mod_6598(clk,rst,matrix_A[6598],matrix_B[198],mul_res1[6598]);
multi_7x28 multi_7x28_mod_6599(clk,rst,matrix_A[6599],matrix_B[199],mul_res1[6599]);
multi_7x28 multi_7x28_mod_6600(clk,rst,matrix_A[6600],matrix_B[0],mul_res1[6600]);
multi_7x28 multi_7x28_mod_6601(clk,rst,matrix_A[6601],matrix_B[1],mul_res1[6601]);
multi_7x28 multi_7x28_mod_6602(clk,rst,matrix_A[6602],matrix_B[2],mul_res1[6602]);
multi_7x28 multi_7x28_mod_6603(clk,rst,matrix_A[6603],matrix_B[3],mul_res1[6603]);
multi_7x28 multi_7x28_mod_6604(clk,rst,matrix_A[6604],matrix_B[4],mul_res1[6604]);
multi_7x28 multi_7x28_mod_6605(clk,rst,matrix_A[6605],matrix_B[5],mul_res1[6605]);
multi_7x28 multi_7x28_mod_6606(clk,rst,matrix_A[6606],matrix_B[6],mul_res1[6606]);
multi_7x28 multi_7x28_mod_6607(clk,rst,matrix_A[6607],matrix_B[7],mul_res1[6607]);
multi_7x28 multi_7x28_mod_6608(clk,rst,matrix_A[6608],matrix_B[8],mul_res1[6608]);
multi_7x28 multi_7x28_mod_6609(clk,rst,matrix_A[6609],matrix_B[9],mul_res1[6609]);
multi_7x28 multi_7x28_mod_6610(clk,rst,matrix_A[6610],matrix_B[10],mul_res1[6610]);
multi_7x28 multi_7x28_mod_6611(clk,rst,matrix_A[6611],matrix_B[11],mul_res1[6611]);
multi_7x28 multi_7x28_mod_6612(clk,rst,matrix_A[6612],matrix_B[12],mul_res1[6612]);
multi_7x28 multi_7x28_mod_6613(clk,rst,matrix_A[6613],matrix_B[13],mul_res1[6613]);
multi_7x28 multi_7x28_mod_6614(clk,rst,matrix_A[6614],matrix_B[14],mul_res1[6614]);
multi_7x28 multi_7x28_mod_6615(clk,rst,matrix_A[6615],matrix_B[15],mul_res1[6615]);
multi_7x28 multi_7x28_mod_6616(clk,rst,matrix_A[6616],matrix_B[16],mul_res1[6616]);
multi_7x28 multi_7x28_mod_6617(clk,rst,matrix_A[6617],matrix_B[17],mul_res1[6617]);
multi_7x28 multi_7x28_mod_6618(clk,rst,matrix_A[6618],matrix_B[18],mul_res1[6618]);
multi_7x28 multi_7x28_mod_6619(clk,rst,matrix_A[6619],matrix_B[19],mul_res1[6619]);
multi_7x28 multi_7x28_mod_6620(clk,rst,matrix_A[6620],matrix_B[20],mul_res1[6620]);
multi_7x28 multi_7x28_mod_6621(clk,rst,matrix_A[6621],matrix_B[21],mul_res1[6621]);
multi_7x28 multi_7x28_mod_6622(clk,rst,matrix_A[6622],matrix_B[22],mul_res1[6622]);
multi_7x28 multi_7x28_mod_6623(clk,rst,matrix_A[6623],matrix_B[23],mul_res1[6623]);
multi_7x28 multi_7x28_mod_6624(clk,rst,matrix_A[6624],matrix_B[24],mul_res1[6624]);
multi_7x28 multi_7x28_mod_6625(clk,rst,matrix_A[6625],matrix_B[25],mul_res1[6625]);
multi_7x28 multi_7x28_mod_6626(clk,rst,matrix_A[6626],matrix_B[26],mul_res1[6626]);
multi_7x28 multi_7x28_mod_6627(clk,rst,matrix_A[6627],matrix_B[27],mul_res1[6627]);
multi_7x28 multi_7x28_mod_6628(clk,rst,matrix_A[6628],matrix_B[28],mul_res1[6628]);
multi_7x28 multi_7x28_mod_6629(clk,rst,matrix_A[6629],matrix_B[29],mul_res1[6629]);
multi_7x28 multi_7x28_mod_6630(clk,rst,matrix_A[6630],matrix_B[30],mul_res1[6630]);
multi_7x28 multi_7x28_mod_6631(clk,rst,matrix_A[6631],matrix_B[31],mul_res1[6631]);
multi_7x28 multi_7x28_mod_6632(clk,rst,matrix_A[6632],matrix_B[32],mul_res1[6632]);
multi_7x28 multi_7x28_mod_6633(clk,rst,matrix_A[6633],matrix_B[33],mul_res1[6633]);
multi_7x28 multi_7x28_mod_6634(clk,rst,matrix_A[6634],matrix_B[34],mul_res1[6634]);
multi_7x28 multi_7x28_mod_6635(clk,rst,matrix_A[6635],matrix_B[35],mul_res1[6635]);
multi_7x28 multi_7x28_mod_6636(clk,rst,matrix_A[6636],matrix_B[36],mul_res1[6636]);
multi_7x28 multi_7x28_mod_6637(clk,rst,matrix_A[6637],matrix_B[37],mul_res1[6637]);
multi_7x28 multi_7x28_mod_6638(clk,rst,matrix_A[6638],matrix_B[38],mul_res1[6638]);
multi_7x28 multi_7x28_mod_6639(clk,rst,matrix_A[6639],matrix_B[39],mul_res1[6639]);
multi_7x28 multi_7x28_mod_6640(clk,rst,matrix_A[6640],matrix_B[40],mul_res1[6640]);
multi_7x28 multi_7x28_mod_6641(clk,rst,matrix_A[6641],matrix_B[41],mul_res1[6641]);
multi_7x28 multi_7x28_mod_6642(clk,rst,matrix_A[6642],matrix_B[42],mul_res1[6642]);
multi_7x28 multi_7x28_mod_6643(clk,rst,matrix_A[6643],matrix_B[43],mul_res1[6643]);
multi_7x28 multi_7x28_mod_6644(clk,rst,matrix_A[6644],matrix_B[44],mul_res1[6644]);
multi_7x28 multi_7x28_mod_6645(clk,rst,matrix_A[6645],matrix_B[45],mul_res1[6645]);
multi_7x28 multi_7x28_mod_6646(clk,rst,matrix_A[6646],matrix_B[46],mul_res1[6646]);
multi_7x28 multi_7x28_mod_6647(clk,rst,matrix_A[6647],matrix_B[47],mul_res1[6647]);
multi_7x28 multi_7x28_mod_6648(clk,rst,matrix_A[6648],matrix_B[48],mul_res1[6648]);
multi_7x28 multi_7x28_mod_6649(clk,rst,matrix_A[6649],matrix_B[49],mul_res1[6649]);
multi_7x28 multi_7x28_mod_6650(clk,rst,matrix_A[6650],matrix_B[50],mul_res1[6650]);
multi_7x28 multi_7x28_mod_6651(clk,rst,matrix_A[6651],matrix_B[51],mul_res1[6651]);
multi_7x28 multi_7x28_mod_6652(clk,rst,matrix_A[6652],matrix_B[52],mul_res1[6652]);
multi_7x28 multi_7x28_mod_6653(clk,rst,matrix_A[6653],matrix_B[53],mul_res1[6653]);
multi_7x28 multi_7x28_mod_6654(clk,rst,matrix_A[6654],matrix_B[54],mul_res1[6654]);
multi_7x28 multi_7x28_mod_6655(clk,rst,matrix_A[6655],matrix_B[55],mul_res1[6655]);
multi_7x28 multi_7x28_mod_6656(clk,rst,matrix_A[6656],matrix_B[56],mul_res1[6656]);
multi_7x28 multi_7x28_mod_6657(clk,rst,matrix_A[6657],matrix_B[57],mul_res1[6657]);
multi_7x28 multi_7x28_mod_6658(clk,rst,matrix_A[6658],matrix_B[58],mul_res1[6658]);
multi_7x28 multi_7x28_mod_6659(clk,rst,matrix_A[6659],matrix_B[59],mul_res1[6659]);
multi_7x28 multi_7x28_mod_6660(clk,rst,matrix_A[6660],matrix_B[60],mul_res1[6660]);
multi_7x28 multi_7x28_mod_6661(clk,rst,matrix_A[6661],matrix_B[61],mul_res1[6661]);
multi_7x28 multi_7x28_mod_6662(clk,rst,matrix_A[6662],matrix_B[62],mul_res1[6662]);
multi_7x28 multi_7x28_mod_6663(clk,rst,matrix_A[6663],matrix_B[63],mul_res1[6663]);
multi_7x28 multi_7x28_mod_6664(clk,rst,matrix_A[6664],matrix_B[64],mul_res1[6664]);
multi_7x28 multi_7x28_mod_6665(clk,rst,matrix_A[6665],matrix_B[65],mul_res1[6665]);
multi_7x28 multi_7x28_mod_6666(clk,rst,matrix_A[6666],matrix_B[66],mul_res1[6666]);
multi_7x28 multi_7x28_mod_6667(clk,rst,matrix_A[6667],matrix_B[67],mul_res1[6667]);
multi_7x28 multi_7x28_mod_6668(clk,rst,matrix_A[6668],matrix_B[68],mul_res1[6668]);
multi_7x28 multi_7x28_mod_6669(clk,rst,matrix_A[6669],matrix_B[69],mul_res1[6669]);
multi_7x28 multi_7x28_mod_6670(clk,rst,matrix_A[6670],matrix_B[70],mul_res1[6670]);
multi_7x28 multi_7x28_mod_6671(clk,rst,matrix_A[6671],matrix_B[71],mul_res1[6671]);
multi_7x28 multi_7x28_mod_6672(clk,rst,matrix_A[6672],matrix_B[72],mul_res1[6672]);
multi_7x28 multi_7x28_mod_6673(clk,rst,matrix_A[6673],matrix_B[73],mul_res1[6673]);
multi_7x28 multi_7x28_mod_6674(clk,rst,matrix_A[6674],matrix_B[74],mul_res1[6674]);
multi_7x28 multi_7x28_mod_6675(clk,rst,matrix_A[6675],matrix_B[75],mul_res1[6675]);
multi_7x28 multi_7x28_mod_6676(clk,rst,matrix_A[6676],matrix_B[76],mul_res1[6676]);
multi_7x28 multi_7x28_mod_6677(clk,rst,matrix_A[6677],matrix_B[77],mul_res1[6677]);
multi_7x28 multi_7x28_mod_6678(clk,rst,matrix_A[6678],matrix_B[78],mul_res1[6678]);
multi_7x28 multi_7x28_mod_6679(clk,rst,matrix_A[6679],matrix_B[79],mul_res1[6679]);
multi_7x28 multi_7x28_mod_6680(clk,rst,matrix_A[6680],matrix_B[80],mul_res1[6680]);
multi_7x28 multi_7x28_mod_6681(clk,rst,matrix_A[6681],matrix_B[81],mul_res1[6681]);
multi_7x28 multi_7x28_mod_6682(clk,rst,matrix_A[6682],matrix_B[82],mul_res1[6682]);
multi_7x28 multi_7x28_mod_6683(clk,rst,matrix_A[6683],matrix_B[83],mul_res1[6683]);
multi_7x28 multi_7x28_mod_6684(clk,rst,matrix_A[6684],matrix_B[84],mul_res1[6684]);
multi_7x28 multi_7x28_mod_6685(clk,rst,matrix_A[6685],matrix_B[85],mul_res1[6685]);
multi_7x28 multi_7x28_mod_6686(clk,rst,matrix_A[6686],matrix_B[86],mul_res1[6686]);
multi_7x28 multi_7x28_mod_6687(clk,rst,matrix_A[6687],matrix_B[87],mul_res1[6687]);
multi_7x28 multi_7x28_mod_6688(clk,rst,matrix_A[6688],matrix_B[88],mul_res1[6688]);
multi_7x28 multi_7x28_mod_6689(clk,rst,matrix_A[6689],matrix_B[89],mul_res1[6689]);
multi_7x28 multi_7x28_mod_6690(clk,rst,matrix_A[6690],matrix_B[90],mul_res1[6690]);
multi_7x28 multi_7x28_mod_6691(clk,rst,matrix_A[6691],matrix_B[91],mul_res1[6691]);
multi_7x28 multi_7x28_mod_6692(clk,rst,matrix_A[6692],matrix_B[92],mul_res1[6692]);
multi_7x28 multi_7x28_mod_6693(clk,rst,matrix_A[6693],matrix_B[93],mul_res1[6693]);
multi_7x28 multi_7x28_mod_6694(clk,rst,matrix_A[6694],matrix_B[94],mul_res1[6694]);
multi_7x28 multi_7x28_mod_6695(clk,rst,matrix_A[6695],matrix_B[95],mul_res1[6695]);
multi_7x28 multi_7x28_mod_6696(clk,rst,matrix_A[6696],matrix_B[96],mul_res1[6696]);
multi_7x28 multi_7x28_mod_6697(clk,rst,matrix_A[6697],matrix_B[97],mul_res1[6697]);
multi_7x28 multi_7x28_mod_6698(clk,rst,matrix_A[6698],matrix_B[98],mul_res1[6698]);
multi_7x28 multi_7x28_mod_6699(clk,rst,matrix_A[6699],matrix_B[99],mul_res1[6699]);
multi_7x28 multi_7x28_mod_6700(clk,rst,matrix_A[6700],matrix_B[100],mul_res1[6700]);
multi_7x28 multi_7x28_mod_6701(clk,rst,matrix_A[6701],matrix_B[101],mul_res1[6701]);
multi_7x28 multi_7x28_mod_6702(clk,rst,matrix_A[6702],matrix_B[102],mul_res1[6702]);
multi_7x28 multi_7x28_mod_6703(clk,rst,matrix_A[6703],matrix_B[103],mul_res1[6703]);
multi_7x28 multi_7x28_mod_6704(clk,rst,matrix_A[6704],matrix_B[104],mul_res1[6704]);
multi_7x28 multi_7x28_mod_6705(clk,rst,matrix_A[6705],matrix_B[105],mul_res1[6705]);
multi_7x28 multi_7x28_mod_6706(clk,rst,matrix_A[6706],matrix_B[106],mul_res1[6706]);
multi_7x28 multi_7x28_mod_6707(clk,rst,matrix_A[6707],matrix_B[107],mul_res1[6707]);
multi_7x28 multi_7x28_mod_6708(clk,rst,matrix_A[6708],matrix_B[108],mul_res1[6708]);
multi_7x28 multi_7x28_mod_6709(clk,rst,matrix_A[6709],matrix_B[109],mul_res1[6709]);
multi_7x28 multi_7x28_mod_6710(clk,rst,matrix_A[6710],matrix_B[110],mul_res1[6710]);
multi_7x28 multi_7x28_mod_6711(clk,rst,matrix_A[6711],matrix_B[111],mul_res1[6711]);
multi_7x28 multi_7x28_mod_6712(clk,rst,matrix_A[6712],matrix_B[112],mul_res1[6712]);
multi_7x28 multi_7x28_mod_6713(clk,rst,matrix_A[6713],matrix_B[113],mul_res1[6713]);
multi_7x28 multi_7x28_mod_6714(clk,rst,matrix_A[6714],matrix_B[114],mul_res1[6714]);
multi_7x28 multi_7x28_mod_6715(clk,rst,matrix_A[6715],matrix_B[115],mul_res1[6715]);
multi_7x28 multi_7x28_mod_6716(clk,rst,matrix_A[6716],matrix_B[116],mul_res1[6716]);
multi_7x28 multi_7x28_mod_6717(clk,rst,matrix_A[6717],matrix_B[117],mul_res1[6717]);
multi_7x28 multi_7x28_mod_6718(clk,rst,matrix_A[6718],matrix_B[118],mul_res1[6718]);
multi_7x28 multi_7x28_mod_6719(clk,rst,matrix_A[6719],matrix_B[119],mul_res1[6719]);
multi_7x28 multi_7x28_mod_6720(clk,rst,matrix_A[6720],matrix_B[120],mul_res1[6720]);
multi_7x28 multi_7x28_mod_6721(clk,rst,matrix_A[6721],matrix_B[121],mul_res1[6721]);
multi_7x28 multi_7x28_mod_6722(clk,rst,matrix_A[6722],matrix_B[122],mul_res1[6722]);
multi_7x28 multi_7x28_mod_6723(clk,rst,matrix_A[6723],matrix_B[123],mul_res1[6723]);
multi_7x28 multi_7x28_mod_6724(clk,rst,matrix_A[6724],matrix_B[124],mul_res1[6724]);
multi_7x28 multi_7x28_mod_6725(clk,rst,matrix_A[6725],matrix_B[125],mul_res1[6725]);
multi_7x28 multi_7x28_mod_6726(clk,rst,matrix_A[6726],matrix_B[126],mul_res1[6726]);
multi_7x28 multi_7x28_mod_6727(clk,rst,matrix_A[6727],matrix_B[127],mul_res1[6727]);
multi_7x28 multi_7x28_mod_6728(clk,rst,matrix_A[6728],matrix_B[128],mul_res1[6728]);
multi_7x28 multi_7x28_mod_6729(clk,rst,matrix_A[6729],matrix_B[129],mul_res1[6729]);
multi_7x28 multi_7x28_mod_6730(clk,rst,matrix_A[6730],matrix_B[130],mul_res1[6730]);
multi_7x28 multi_7x28_mod_6731(clk,rst,matrix_A[6731],matrix_B[131],mul_res1[6731]);
multi_7x28 multi_7x28_mod_6732(clk,rst,matrix_A[6732],matrix_B[132],mul_res1[6732]);
multi_7x28 multi_7x28_mod_6733(clk,rst,matrix_A[6733],matrix_B[133],mul_res1[6733]);
multi_7x28 multi_7x28_mod_6734(clk,rst,matrix_A[6734],matrix_B[134],mul_res1[6734]);
multi_7x28 multi_7x28_mod_6735(clk,rst,matrix_A[6735],matrix_B[135],mul_res1[6735]);
multi_7x28 multi_7x28_mod_6736(clk,rst,matrix_A[6736],matrix_B[136],mul_res1[6736]);
multi_7x28 multi_7x28_mod_6737(clk,rst,matrix_A[6737],matrix_B[137],mul_res1[6737]);
multi_7x28 multi_7x28_mod_6738(clk,rst,matrix_A[6738],matrix_B[138],mul_res1[6738]);
multi_7x28 multi_7x28_mod_6739(clk,rst,matrix_A[6739],matrix_B[139],mul_res1[6739]);
multi_7x28 multi_7x28_mod_6740(clk,rst,matrix_A[6740],matrix_B[140],mul_res1[6740]);
multi_7x28 multi_7x28_mod_6741(clk,rst,matrix_A[6741],matrix_B[141],mul_res1[6741]);
multi_7x28 multi_7x28_mod_6742(clk,rst,matrix_A[6742],matrix_B[142],mul_res1[6742]);
multi_7x28 multi_7x28_mod_6743(clk,rst,matrix_A[6743],matrix_B[143],mul_res1[6743]);
multi_7x28 multi_7x28_mod_6744(clk,rst,matrix_A[6744],matrix_B[144],mul_res1[6744]);
multi_7x28 multi_7x28_mod_6745(clk,rst,matrix_A[6745],matrix_B[145],mul_res1[6745]);
multi_7x28 multi_7x28_mod_6746(clk,rst,matrix_A[6746],matrix_B[146],mul_res1[6746]);
multi_7x28 multi_7x28_mod_6747(clk,rst,matrix_A[6747],matrix_B[147],mul_res1[6747]);
multi_7x28 multi_7x28_mod_6748(clk,rst,matrix_A[6748],matrix_B[148],mul_res1[6748]);
multi_7x28 multi_7x28_mod_6749(clk,rst,matrix_A[6749],matrix_B[149],mul_res1[6749]);
multi_7x28 multi_7x28_mod_6750(clk,rst,matrix_A[6750],matrix_B[150],mul_res1[6750]);
multi_7x28 multi_7x28_mod_6751(clk,rst,matrix_A[6751],matrix_B[151],mul_res1[6751]);
multi_7x28 multi_7x28_mod_6752(clk,rst,matrix_A[6752],matrix_B[152],mul_res1[6752]);
multi_7x28 multi_7x28_mod_6753(clk,rst,matrix_A[6753],matrix_B[153],mul_res1[6753]);
multi_7x28 multi_7x28_mod_6754(clk,rst,matrix_A[6754],matrix_B[154],mul_res1[6754]);
multi_7x28 multi_7x28_mod_6755(clk,rst,matrix_A[6755],matrix_B[155],mul_res1[6755]);
multi_7x28 multi_7x28_mod_6756(clk,rst,matrix_A[6756],matrix_B[156],mul_res1[6756]);
multi_7x28 multi_7x28_mod_6757(clk,rst,matrix_A[6757],matrix_B[157],mul_res1[6757]);
multi_7x28 multi_7x28_mod_6758(clk,rst,matrix_A[6758],matrix_B[158],mul_res1[6758]);
multi_7x28 multi_7x28_mod_6759(clk,rst,matrix_A[6759],matrix_B[159],mul_res1[6759]);
multi_7x28 multi_7x28_mod_6760(clk,rst,matrix_A[6760],matrix_B[160],mul_res1[6760]);
multi_7x28 multi_7x28_mod_6761(clk,rst,matrix_A[6761],matrix_B[161],mul_res1[6761]);
multi_7x28 multi_7x28_mod_6762(clk,rst,matrix_A[6762],matrix_B[162],mul_res1[6762]);
multi_7x28 multi_7x28_mod_6763(clk,rst,matrix_A[6763],matrix_B[163],mul_res1[6763]);
multi_7x28 multi_7x28_mod_6764(clk,rst,matrix_A[6764],matrix_B[164],mul_res1[6764]);
multi_7x28 multi_7x28_mod_6765(clk,rst,matrix_A[6765],matrix_B[165],mul_res1[6765]);
multi_7x28 multi_7x28_mod_6766(clk,rst,matrix_A[6766],matrix_B[166],mul_res1[6766]);
multi_7x28 multi_7x28_mod_6767(clk,rst,matrix_A[6767],matrix_B[167],mul_res1[6767]);
multi_7x28 multi_7x28_mod_6768(clk,rst,matrix_A[6768],matrix_B[168],mul_res1[6768]);
multi_7x28 multi_7x28_mod_6769(clk,rst,matrix_A[6769],matrix_B[169],mul_res1[6769]);
multi_7x28 multi_7x28_mod_6770(clk,rst,matrix_A[6770],matrix_B[170],mul_res1[6770]);
multi_7x28 multi_7x28_mod_6771(clk,rst,matrix_A[6771],matrix_B[171],mul_res1[6771]);
multi_7x28 multi_7x28_mod_6772(clk,rst,matrix_A[6772],matrix_B[172],mul_res1[6772]);
multi_7x28 multi_7x28_mod_6773(clk,rst,matrix_A[6773],matrix_B[173],mul_res1[6773]);
multi_7x28 multi_7x28_mod_6774(clk,rst,matrix_A[6774],matrix_B[174],mul_res1[6774]);
multi_7x28 multi_7x28_mod_6775(clk,rst,matrix_A[6775],matrix_B[175],mul_res1[6775]);
multi_7x28 multi_7x28_mod_6776(clk,rst,matrix_A[6776],matrix_B[176],mul_res1[6776]);
multi_7x28 multi_7x28_mod_6777(clk,rst,matrix_A[6777],matrix_B[177],mul_res1[6777]);
multi_7x28 multi_7x28_mod_6778(clk,rst,matrix_A[6778],matrix_B[178],mul_res1[6778]);
multi_7x28 multi_7x28_mod_6779(clk,rst,matrix_A[6779],matrix_B[179],mul_res1[6779]);
multi_7x28 multi_7x28_mod_6780(clk,rst,matrix_A[6780],matrix_B[180],mul_res1[6780]);
multi_7x28 multi_7x28_mod_6781(clk,rst,matrix_A[6781],matrix_B[181],mul_res1[6781]);
multi_7x28 multi_7x28_mod_6782(clk,rst,matrix_A[6782],matrix_B[182],mul_res1[6782]);
multi_7x28 multi_7x28_mod_6783(clk,rst,matrix_A[6783],matrix_B[183],mul_res1[6783]);
multi_7x28 multi_7x28_mod_6784(clk,rst,matrix_A[6784],matrix_B[184],mul_res1[6784]);
multi_7x28 multi_7x28_mod_6785(clk,rst,matrix_A[6785],matrix_B[185],mul_res1[6785]);
multi_7x28 multi_7x28_mod_6786(clk,rst,matrix_A[6786],matrix_B[186],mul_res1[6786]);
multi_7x28 multi_7x28_mod_6787(clk,rst,matrix_A[6787],matrix_B[187],mul_res1[6787]);
multi_7x28 multi_7x28_mod_6788(clk,rst,matrix_A[6788],matrix_B[188],mul_res1[6788]);
multi_7x28 multi_7x28_mod_6789(clk,rst,matrix_A[6789],matrix_B[189],mul_res1[6789]);
multi_7x28 multi_7x28_mod_6790(clk,rst,matrix_A[6790],matrix_B[190],mul_res1[6790]);
multi_7x28 multi_7x28_mod_6791(clk,rst,matrix_A[6791],matrix_B[191],mul_res1[6791]);
multi_7x28 multi_7x28_mod_6792(clk,rst,matrix_A[6792],matrix_B[192],mul_res1[6792]);
multi_7x28 multi_7x28_mod_6793(clk,rst,matrix_A[6793],matrix_B[193],mul_res1[6793]);
multi_7x28 multi_7x28_mod_6794(clk,rst,matrix_A[6794],matrix_B[194],mul_res1[6794]);
multi_7x28 multi_7x28_mod_6795(clk,rst,matrix_A[6795],matrix_B[195],mul_res1[6795]);
multi_7x28 multi_7x28_mod_6796(clk,rst,matrix_A[6796],matrix_B[196],mul_res1[6796]);
multi_7x28 multi_7x28_mod_6797(clk,rst,matrix_A[6797],matrix_B[197],mul_res1[6797]);
multi_7x28 multi_7x28_mod_6798(clk,rst,matrix_A[6798],matrix_B[198],mul_res1[6798]);
multi_7x28 multi_7x28_mod_6799(clk,rst,matrix_A[6799],matrix_B[199],mul_res1[6799]);
multi_7x28 multi_7x28_mod_6800(clk,rst,matrix_A[6800],matrix_B[0],mul_res1[6800]);
multi_7x28 multi_7x28_mod_6801(clk,rst,matrix_A[6801],matrix_B[1],mul_res1[6801]);
multi_7x28 multi_7x28_mod_6802(clk,rst,matrix_A[6802],matrix_B[2],mul_res1[6802]);
multi_7x28 multi_7x28_mod_6803(clk,rst,matrix_A[6803],matrix_B[3],mul_res1[6803]);
multi_7x28 multi_7x28_mod_6804(clk,rst,matrix_A[6804],matrix_B[4],mul_res1[6804]);
multi_7x28 multi_7x28_mod_6805(clk,rst,matrix_A[6805],matrix_B[5],mul_res1[6805]);
multi_7x28 multi_7x28_mod_6806(clk,rst,matrix_A[6806],matrix_B[6],mul_res1[6806]);
multi_7x28 multi_7x28_mod_6807(clk,rst,matrix_A[6807],matrix_B[7],mul_res1[6807]);
multi_7x28 multi_7x28_mod_6808(clk,rst,matrix_A[6808],matrix_B[8],mul_res1[6808]);
multi_7x28 multi_7x28_mod_6809(clk,rst,matrix_A[6809],matrix_B[9],mul_res1[6809]);
multi_7x28 multi_7x28_mod_6810(clk,rst,matrix_A[6810],matrix_B[10],mul_res1[6810]);
multi_7x28 multi_7x28_mod_6811(clk,rst,matrix_A[6811],matrix_B[11],mul_res1[6811]);
multi_7x28 multi_7x28_mod_6812(clk,rst,matrix_A[6812],matrix_B[12],mul_res1[6812]);
multi_7x28 multi_7x28_mod_6813(clk,rst,matrix_A[6813],matrix_B[13],mul_res1[6813]);
multi_7x28 multi_7x28_mod_6814(clk,rst,matrix_A[6814],matrix_B[14],mul_res1[6814]);
multi_7x28 multi_7x28_mod_6815(clk,rst,matrix_A[6815],matrix_B[15],mul_res1[6815]);
multi_7x28 multi_7x28_mod_6816(clk,rst,matrix_A[6816],matrix_B[16],mul_res1[6816]);
multi_7x28 multi_7x28_mod_6817(clk,rst,matrix_A[6817],matrix_B[17],mul_res1[6817]);
multi_7x28 multi_7x28_mod_6818(clk,rst,matrix_A[6818],matrix_B[18],mul_res1[6818]);
multi_7x28 multi_7x28_mod_6819(clk,rst,matrix_A[6819],matrix_B[19],mul_res1[6819]);
multi_7x28 multi_7x28_mod_6820(clk,rst,matrix_A[6820],matrix_B[20],mul_res1[6820]);
multi_7x28 multi_7x28_mod_6821(clk,rst,matrix_A[6821],matrix_B[21],mul_res1[6821]);
multi_7x28 multi_7x28_mod_6822(clk,rst,matrix_A[6822],matrix_B[22],mul_res1[6822]);
multi_7x28 multi_7x28_mod_6823(clk,rst,matrix_A[6823],matrix_B[23],mul_res1[6823]);
multi_7x28 multi_7x28_mod_6824(clk,rst,matrix_A[6824],matrix_B[24],mul_res1[6824]);
multi_7x28 multi_7x28_mod_6825(clk,rst,matrix_A[6825],matrix_B[25],mul_res1[6825]);
multi_7x28 multi_7x28_mod_6826(clk,rst,matrix_A[6826],matrix_B[26],mul_res1[6826]);
multi_7x28 multi_7x28_mod_6827(clk,rst,matrix_A[6827],matrix_B[27],mul_res1[6827]);
multi_7x28 multi_7x28_mod_6828(clk,rst,matrix_A[6828],matrix_B[28],mul_res1[6828]);
multi_7x28 multi_7x28_mod_6829(clk,rst,matrix_A[6829],matrix_B[29],mul_res1[6829]);
multi_7x28 multi_7x28_mod_6830(clk,rst,matrix_A[6830],matrix_B[30],mul_res1[6830]);
multi_7x28 multi_7x28_mod_6831(clk,rst,matrix_A[6831],matrix_B[31],mul_res1[6831]);
multi_7x28 multi_7x28_mod_6832(clk,rst,matrix_A[6832],matrix_B[32],mul_res1[6832]);
multi_7x28 multi_7x28_mod_6833(clk,rst,matrix_A[6833],matrix_B[33],mul_res1[6833]);
multi_7x28 multi_7x28_mod_6834(clk,rst,matrix_A[6834],matrix_B[34],mul_res1[6834]);
multi_7x28 multi_7x28_mod_6835(clk,rst,matrix_A[6835],matrix_B[35],mul_res1[6835]);
multi_7x28 multi_7x28_mod_6836(clk,rst,matrix_A[6836],matrix_B[36],mul_res1[6836]);
multi_7x28 multi_7x28_mod_6837(clk,rst,matrix_A[6837],matrix_B[37],mul_res1[6837]);
multi_7x28 multi_7x28_mod_6838(clk,rst,matrix_A[6838],matrix_B[38],mul_res1[6838]);
multi_7x28 multi_7x28_mod_6839(clk,rst,matrix_A[6839],matrix_B[39],mul_res1[6839]);
multi_7x28 multi_7x28_mod_6840(clk,rst,matrix_A[6840],matrix_B[40],mul_res1[6840]);
multi_7x28 multi_7x28_mod_6841(clk,rst,matrix_A[6841],matrix_B[41],mul_res1[6841]);
multi_7x28 multi_7x28_mod_6842(clk,rst,matrix_A[6842],matrix_B[42],mul_res1[6842]);
multi_7x28 multi_7x28_mod_6843(clk,rst,matrix_A[6843],matrix_B[43],mul_res1[6843]);
multi_7x28 multi_7x28_mod_6844(clk,rst,matrix_A[6844],matrix_B[44],mul_res1[6844]);
multi_7x28 multi_7x28_mod_6845(clk,rst,matrix_A[6845],matrix_B[45],mul_res1[6845]);
multi_7x28 multi_7x28_mod_6846(clk,rst,matrix_A[6846],matrix_B[46],mul_res1[6846]);
multi_7x28 multi_7x28_mod_6847(clk,rst,matrix_A[6847],matrix_B[47],mul_res1[6847]);
multi_7x28 multi_7x28_mod_6848(clk,rst,matrix_A[6848],matrix_B[48],mul_res1[6848]);
multi_7x28 multi_7x28_mod_6849(clk,rst,matrix_A[6849],matrix_B[49],mul_res1[6849]);
multi_7x28 multi_7x28_mod_6850(clk,rst,matrix_A[6850],matrix_B[50],mul_res1[6850]);
multi_7x28 multi_7x28_mod_6851(clk,rst,matrix_A[6851],matrix_B[51],mul_res1[6851]);
multi_7x28 multi_7x28_mod_6852(clk,rst,matrix_A[6852],matrix_B[52],mul_res1[6852]);
multi_7x28 multi_7x28_mod_6853(clk,rst,matrix_A[6853],matrix_B[53],mul_res1[6853]);
multi_7x28 multi_7x28_mod_6854(clk,rst,matrix_A[6854],matrix_B[54],mul_res1[6854]);
multi_7x28 multi_7x28_mod_6855(clk,rst,matrix_A[6855],matrix_B[55],mul_res1[6855]);
multi_7x28 multi_7x28_mod_6856(clk,rst,matrix_A[6856],matrix_B[56],mul_res1[6856]);
multi_7x28 multi_7x28_mod_6857(clk,rst,matrix_A[6857],matrix_B[57],mul_res1[6857]);
multi_7x28 multi_7x28_mod_6858(clk,rst,matrix_A[6858],matrix_B[58],mul_res1[6858]);
multi_7x28 multi_7x28_mod_6859(clk,rst,matrix_A[6859],matrix_B[59],mul_res1[6859]);
multi_7x28 multi_7x28_mod_6860(clk,rst,matrix_A[6860],matrix_B[60],mul_res1[6860]);
multi_7x28 multi_7x28_mod_6861(clk,rst,matrix_A[6861],matrix_B[61],mul_res1[6861]);
multi_7x28 multi_7x28_mod_6862(clk,rst,matrix_A[6862],matrix_B[62],mul_res1[6862]);
multi_7x28 multi_7x28_mod_6863(clk,rst,matrix_A[6863],matrix_B[63],mul_res1[6863]);
multi_7x28 multi_7x28_mod_6864(clk,rst,matrix_A[6864],matrix_B[64],mul_res1[6864]);
multi_7x28 multi_7x28_mod_6865(clk,rst,matrix_A[6865],matrix_B[65],mul_res1[6865]);
multi_7x28 multi_7x28_mod_6866(clk,rst,matrix_A[6866],matrix_B[66],mul_res1[6866]);
multi_7x28 multi_7x28_mod_6867(clk,rst,matrix_A[6867],matrix_B[67],mul_res1[6867]);
multi_7x28 multi_7x28_mod_6868(clk,rst,matrix_A[6868],matrix_B[68],mul_res1[6868]);
multi_7x28 multi_7x28_mod_6869(clk,rst,matrix_A[6869],matrix_B[69],mul_res1[6869]);
multi_7x28 multi_7x28_mod_6870(clk,rst,matrix_A[6870],matrix_B[70],mul_res1[6870]);
multi_7x28 multi_7x28_mod_6871(clk,rst,matrix_A[6871],matrix_B[71],mul_res1[6871]);
multi_7x28 multi_7x28_mod_6872(clk,rst,matrix_A[6872],matrix_B[72],mul_res1[6872]);
multi_7x28 multi_7x28_mod_6873(clk,rst,matrix_A[6873],matrix_B[73],mul_res1[6873]);
multi_7x28 multi_7x28_mod_6874(clk,rst,matrix_A[6874],matrix_B[74],mul_res1[6874]);
multi_7x28 multi_7x28_mod_6875(clk,rst,matrix_A[6875],matrix_B[75],mul_res1[6875]);
multi_7x28 multi_7x28_mod_6876(clk,rst,matrix_A[6876],matrix_B[76],mul_res1[6876]);
multi_7x28 multi_7x28_mod_6877(clk,rst,matrix_A[6877],matrix_B[77],mul_res1[6877]);
multi_7x28 multi_7x28_mod_6878(clk,rst,matrix_A[6878],matrix_B[78],mul_res1[6878]);
multi_7x28 multi_7x28_mod_6879(clk,rst,matrix_A[6879],matrix_B[79],mul_res1[6879]);
multi_7x28 multi_7x28_mod_6880(clk,rst,matrix_A[6880],matrix_B[80],mul_res1[6880]);
multi_7x28 multi_7x28_mod_6881(clk,rst,matrix_A[6881],matrix_B[81],mul_res1[6881]);
multi_7x28 multi_7x28_mod_6882(clk,rst,matrix_A[6882],matrix_B[82],mul_res1[6882]);
multi_7x28 multi_7x28_mod_6883(clk,rst,matrix_A[6883],matrix_B[83],mul_res1[6883]);
multi_7x28 multi_7x28_mod_6884(clk,rst,matrix_A[6884],matrix_B[84],mul_res1[6884]);
multi_7x28 multi_7x28_mod_6885(clk,rst,matrix_A[6885],matrix_B[85],mul_res1[6885]);
multi_7x28 multi_7x28_mod_6886(clk,rst,matrix_A[6886],matrix_B[86],mul_res1[6886]);
multi_7x28 multi_7x28_mod_6887(clk,rst,matrix_A[6887],matrix_B[87],mul_res1[6887]);
multi_7x28 multi_7x28_mod_6888(clk,rst,matrix_A[6888],matrix_B[88],mul_res1[6888]);
multi_7x28 multi_7x28_mod_6889(clk,rst,matrix_A[6889],matrix_B[89],mul_res1[6889]);
multi_7x28 multi_7x28_mod_6890(clk,rst,matrix_A[6890],matrix_B[90],mul_res1[6890]);
multi_7x28 multi_7x28_mod_6891(clk,rst,matrix_A[6891],matrix_B[91],mul_res1[6891]);
multi_7x28 multi_7x28_mod_6892(clk,rst,matrix_A[6892],matrix_B[92],mul_res1[6892]);
multi_7x28 multi_7x28_mod_6893(clk,rst,matrix_A[6893],matrix_B[93],mul_res1[6893]);
multi_7x28 multi_7x28_mod_6894(clk,rst,matrix_A[6894],matrix_B[94],mul_res1[6894]);
multi_7x28 multi_7x28_mod_6895(clk,rst,matrix_A[6895],matrix_B[95],mul_res1[6895]);
multi_7x28 multi_7x28_mod_6896(clk,rst,matrix_A[6896],matrix_B[96],mul_res1[6896]);
multi_7x28 multi_7x28_mod_6897(clk,rst,matrix_A[6897],matrix_B[97],mul_res1[6897]);
multi_7x28 multi_7x28_mod_6898(clk,rst,matrix_A[6898],matrix_B[98],mul_res1[6898]);
multi_7x28 multi_7x28_mod_6899(clk,rst,matrix_A[6899],matrix_B[99],mul_res1[6899]);
multi_7x28 multi_7x28_mod_6900(clk,rst,matrix_A[6900],matrix_B[100],mul_res1[6900]);
multi_7x28 multi_7x28_mod_6901(clk,rst,matrix_A[6901],matrix_B[101],mul_res1[6901]);
multi_7x28 multi_7x28_mod_6902(clk,rst,matrix_A[6902],matrix_B[102],mul_res1[6902]);
multi_7x28 multi_7x28_mod_6903(clk,rst,matrix_A[6903],matrix_B[103],mul_res1[6903]);
multi_7x28 multi_7x28_mod_6904(clk,rst,matrix_A[6904],matrix_B[104],mul_res1[6904]);
multi_7x28 multi_7x28_mod_6905(clk,rst,matrix_A[6905],matrix_B[105],mul_res1[6905]);
multi_7x28 multi_7x28_mod_6906(clk,rst,matrix_A[6906],matrix_B[106],mul_res1[6906]);
multi_7x28 multi_7x28_mod_6907(clk,rst,matrix_A[6907],matrix_B[107],mul_res1[6907]);
multi_7x28 multi_7x28_mod_6908(clk,rst,matrix_A[6908],matrix_B[108],mul_res1[6908]);
multi_7x28 multi_7x28_mod_6909(clk,rst,matrix_A[6909],matrix_B[109],mul_res1[6909]);
multi_7x28 multi_7x28_mod_6910(clk,rst,matrix_A[6910],matrix_B[110],mul_res1[6910]);
multi_7x28 multi_7x28_mod_6911(clk,rst,matrix_A[6911],matrix_B[111],mul_res1[6911]);
multi_7x28 multi_7x28_mod_6912(clk,rst,matrix_A[6912],matrix_B[112],mul_res1[6912]);
multi_7x28 multi_7x28_mod_6913(clk,rst,matrix_A[6913],matrix_B[113],mul_res1[6913]);
multi_7x28 multi_7x28_mod_6914(clk,rst,matrix_A[6914],matrix_B[114],mul_res1[6914]);
multi_7x28 multi_7x28_mod_6915(clk,rst,matrix_A[6915],matrix_B[115],mul_res1[6915]);
multi_7x28 multi_7x28_mod_6916(clk,rst,matrix_A[6916],matrix_B[116],mul_res1[6916]);
multi_7x28 multi_7x28_mod_6917(clk,rst,matrix_A[6917],matrix_B[117],mul_res1[6917]);
multi_7x28 multi_7x28_mod_6918(clk,rst,matrix_A[6918],matrix_B[118],mul_res1[6918]);
multi_7x28 multi_7x28_mod_6919(clk,rst,matrix_A[6919],matrix_B[119],mul_res1[6919]);
multi_7x28 multi_7x28_mod_6920(clk,rst,matrix_A[6920],matrix_B[120],mul_res1[6920]);
multi_7x28 multi_7x28_mod_6921(clk,rst,matrix_A[6921],matrix_B[121],mul_res1[6921]);
multi_7x28 multi_7x28_mod_6922(clk,rst,matrix_A[6922],matrix_B[122],mul_res1[6922]);
multi_7x28 multi_7x28_mod_6923(clk,rst,matrix_A[6923],matrix_B[123],mul_res1[6923]);
multi_7x28 multi_7x28_mod_6924(clk,rst,matrix_A[6924],matrix_B[124],mul_res1[6924]);
multi_7x28 multi_7x28_mod_6925(clk,rst,matrix_A[6925],matrix_B[125],mul_res1[6925]);
multi_7x28 multi_7x28_mod_6926(clk,rst,matrix_A[6926],matrix_B[126],mul_res1[6926]);
multi_7x28 multi_7x28_mod_6927(clk,rst,matrix_A[6927],matrix_B[127],mul_res1[6927]);
multi_7x28 multi_7x28_mod_6928(clk,rst,matrix_A[6928],matrix_B[128],mul_res1[6928]);
multi_7x28 multi_7x28_mod_6929(clk,rst,matrix_A[6929],matrix_B[129],mul_res1[6929]);
multi_7x28 multi_7x28_mod_6930(clk,rst,matrix_A[6930],matrix_B[130],mul_res1[6930]);
multi_7x28 multi_7x28_mod_6931(clk,rst,matrix_A[6931],matrix_B[131],mul_res1[6931]);
multi_7x28 multi_7x28_mod_6932(clk,rst,matrix_A[6932],matrix_B[132],mul_res1[6932]);
multi_7x28 multi_7x28_mod_6933(clk,rst,matrix_A[6933],matrix_B[133],mul_res1[6933]);
multi_7x28 multi_7x28_mod_6934(clk,rst,matrix_A[6934],matrix_B[134],mul_res1[6934]);
multi_7x28 multi_7x28_mod_6935(clk,rst,matrix_A[6935],matrix_B[135],mul_res1[6935]);
multi_7x28 multi_7x28_mod_6936(clk,rst,matrix_A[6936],matrix_B[136],mul_res1[6936]);
multi_7x28 multi_7x28_mod_6937(clk,rst,matrix_A[6937],matrix_B[137],mul_res1[6937]);
multi_7x28 multi_7x28_mod_6938(clk,rst,matrix_A[6938],matrix_B[138],mul_res1[6938]);
multi_7x28 multi_7x28_mod_6939(clk,rst,matrix_A[6939],matrix_B[139],mul_res1[6939]);
multi_7x28 multi_7x28_mod_6940(clk,rst,matrix_A[6940],matrix_B[140],mul_res1[6940]);
multi_7x28 multi_7x28_mod_6941(clk,rst,matrix_A[6941],matrix_B[141],mul_res1[6941]);
multi_7x28 multi_7x28_mod_6942(clk,rst,matrix_A[6942],matrix_B[142],mul_res1[6942]);
multi_7x28 multi_7x28_mod_6943(clk,rst,matrix_A[6943],matrix_B[143],mul_res1[6943]);
multi_7x28 multi_7x28_mod_6944(clk,rst,matrix_A[6944],matrix_B[144],mul_res1[6944]);
multi_7x28 multi_7x28_mod_6945(clk,rst,matrix_A[6945],matrix_B[145],mul_res1[6945]);
multi_7x28 multi_7x28_mod_6946(clk,rst,matrix_A[6946],matrix_B[146],mul_res1[6946]);
multi_7x28 multi_7x28_mod_6947(clk,rst,matrix_A[6947],matrix_B[147],mul_res1[6947]);
multi_7x28 multi_7x28_mod_6948(clk,rst,matrix_A[6948],matrix_B[148],mul_res1[6948]);
multi_7x28 multi_7x28_mod_6949(clk,rst,matrix_A[6949],matrix_B[149],mul_res1[6949]);
multi_7x28 multi_7x28_mod_6950(clk,rst,matrix_A[6950],matrix_B[150],mul_res1[6950]);
multi_7x28 multi_7x28_mod_6951(clk,rst,matrix_A[6951],matrix_B[151],mul_res1[6951]);
multi_7x28 multi_7x28_mod_6952(clk,rst,matrix_A[6952],matrix_B[152],mul_res1[6952]);
multi_7x28 multi_7x28_mod_6953(clk,rst,matrix_A[6953],matrix_B[153],mul_res1[6953]);
multi_7x28 multi_7x28_mod_6954(clk,rst,matrix_A[6954],matrix_B[154],mul_res1[6954]);
multi_7x28 multi_7x28_mod_6955(clk,rst,matrix_A[6955],matrix_B[155],mul_res1[6955]);
multi_7x28 multi_7x28_mod_6956(clk,rst,matrix_A[6956],matrix_B[156],mul_res1[6956]);
multi_7x28 multi_7x28_mod_6957(clk,rst,matrix_A[6957],matrix_B[157],mul_res1[6957]);
multi_7x28 multi_7x28_mod_6958(clk,rst,matrix_A[6958],matrix_B[158],mul_res1[6958]);
multi_7x28 multi_7x28_mod_6959(clk,rst,matrix_A[6959],matrix_B[159],mul_res1[6959]);
multi_7x28 multi_7x28_mod_6960(clk,rst,matrix_A[6960],matrix_B[160],mul_res1[6960]);
multi_7x28 multi_7x28_mod_6961(clk,rst,matrix_A[6961],matrix_B[161],mul_res1[6961]);
multi_7x28 multi_7x28_mod_6962(clk,rst,matrix_A[6962],matrix_B[162],mul_res1[6962]);
multi_7x28 multi_7x28_mod_6963(clk,rst,matrix_A[6963],matrix_B[163],mul_res1[6963]);
multi_7x28 multi_7x28_mod_6964(clk,rst,matrix_A[6964],matrix_B[164],mul_res1[6964]);
multi_7x28 multi_7x28_mod_6965(clk,rst,matrix_A[6965],matrix_B[165],mul_res1[6965]);
multi_7x28 multi_7x28_mod_6966(clk,rst,matrix_A[6966],matrix_B[166],mul_res1[6966]);
multi_7x28 multi_7x28_mod_6967(clk,rst,matrix_A[6967],matrix_B[167],mul_res1[6967]);
multi_7x28 multi_7x28_mod_6968(clk,rst,matrix_A[6968],matrix_B[168],mul_res1[6968]);
multi_7x28 multi_7x28_mod_6969(clk,rst,matrix_A[6969],matrix_B[169],mul_res1[6969]);
multi_7x28 multi_7x28_mod_6970(clk,rst,matrix_A[6970],matrix_B[170],mul_res1[6970]);
multi_7x28 multi_7x28_mod_6971(clk,rst,matrix_A[6971],matrix_B[171],mul_res1[6971]);
multi_7x28 multi_7x28_mod_6972(clk,rst,matrix_A[6972],matrix_B[172],mul_res1[6972]);
multi_7x28 multi_7x28_mod_6973(clk,rst,matrix_A[6973],matrix_B[173],mul_res1[6973]);
multi_7x28 multi_7x28_mod_6974(clk,rst,matrix_A[6974],matrix_B[174],mul_res1[6974]);
multi_7x28 multi_7x28_mod_6975(clk,rst,matrix_A[6975],matrix_B[175],mul_res1[6975]);
multi_7x28 multi_7x28_mod_6976(clk,rst,matrix_A[6976],matrix_B[176],mul_res1[6976]);
multi_7x28 multi_7x28_mod_6977(clk,rst,matrix_A[6977],matrix_B[177],mul_res1[6977]);
multi_7x28 multi_7x28_mod_6978(clk,rst,matrix_A[6978],matrix_B[178],mul_res1[6978]);
multi_7x28 multi_7x28_mod_6979(clk,rst,matrix_A[6979],matrix_B[179],mul_res1[6979]);
multi_7x28 multi_7x28_mod_6980(clk,rst,matrix_A[6980],matrix_B[180],mul_res1[6980]);
multi_7x28 multi_7x28_mod_6981(clk,rst,matrix_A[6981],matrix_B[181],mul_res1[6981]);
multi_7x28 multi_7x28_mod_6982(clk,rst,matrix_A[6982],matrix_B[182],mul_res1[6982]);
multi_7x28 multi_7x28_mod_6983(clk,rst,matrix_A[6983],matrix_B[183],mul_res1[6983]);
multi_7x28 multi_7x28_mod_6984(clk,rst,matrix_A[6984],matrix_B[184],mul_res1[6984]);
multi_7x28 multi_7x28_mod_6985(clk,rst,matrix_A[6985],matrix_B[185],mul_res1[6985]);
multi_7x28 multi_7x28_mod_6986(clk,rst,matrix_A[6986],matrix_B[186],mul_res1[6986]);
multi_7x28 multi_7x28_mod_6987(clk,rst,matrix_A[6987],matrix_B[187],mul_res1[6987]);
multi_7x28 multi_7x28_mod_6988(clk,rst,matrix_A[6988],matrix_B[188],mul_res1[6988]);
multi_7x28 multi_7x28_mod_6989(clk,rst,matrix_A[6989],matrix_B[189],mul_res1[6989]);
multi_7x28 multi_7x28_mod_6990(clk,rst,matrix_A[6990],matrix_B[190],mul_res1[6990]);
multi_7x28 multi_7x28_mod_6991(clk,rst,matrix_A[6991],matrix_B[191],mul_res1[6991]);
multi_7x28 multi_7x28_mod_6992(clk,rst,matrix_A[6992],matrix_B[192],mul_res1[6992]);
multi_7x28 multi_7x28_mod_6993(clk,rst,matrix_A[6993],matrix_B[193],mul_res1[6993]);
multi_7x28 multi_7x28_mod_6994(clk,rst,matrix_A[6994],matrix_B[194],mul_res1[6994]);
multi_7x28 multi_7x28_mod_6995(clk,rst,matrix_A[6995],matrix_B[195],mul_res1[6995]);
multi_7x28 multi_7x28_mod_6996(clk,rst,matrix_A[6996],matrix_B[196],mul_res1[6996]);
multi_7x28 multi_7x28_mod_6997(clk,rst,matrix_A[6997],matrix_B[197],mul_res1[6997]);
multi_7x28 multi_7x28_mod_6998(clk,rst,matrix_A[6998],matrix_B[198],mul_res1[6998]);
multi_7x28 multi_7x28_mod_6999(clk,rst,matrix_A[6999],matrix_B[199],mul_res1[6999]);
multi_7x28 multi_7x28_mod_7000(clk,rst,matrix_A[7000],matrix_B[0],mul_res1[7000]);
multi_7x28 multi_7x28_mod_7001(clk,rst,matrix_A[7001],matrix_B[1],mul_res1[7001]);
multi_7x28 multi_7x28_mod_7002(clk,rst,matrix_A[7002],matrix_B[2],mul_res1[7002]);
multi_7x28 multi_7x28_mod_7003(clk,rst,matrix_A[7003],matrix_B[3],mul_res1[7003]);
multi_7x28 multi_7x28_mod_7004(clk,rst,matrix_A[7004],matrix_B[4],mul_res1[7004]);
multi_7x28 multi_7x28_mod_7005(clk,rst,matrix_A[7005],matrix_B[5],mul_res1[7005]);
multi_7x28 multi_7x28_mod_7006(clk,rst,matrix_A[7006],matrix_B[6],mul_res1[7006]);
multi_7x28 multi_7x28_mod_7007(clk,rst,matrix_A[7007],matrix_B[7],mul_res1[7007]);
multi_7x28 multi_7x28_mod_7008(clk,rst,matrix_A[7008],matrix_B[8],mul_res1[7008]);
multi_7x28 multi_7x28_mod_7009(clk,rst,matrix_A[7009],matrix_B[9],mul_res1[7009]);
multi_7x28 multi_7x28_mod_7010(clk,rst,matrix_A[7010],matrix_B[10],mul_res1[7010]);
multi_7x28 multi_7x28_mod_7011(clk,rst,matrix_A[7011],matrix_B[11],mul_res1[7011]);
multi_7x28 multi_7x28_mod_7012(clk,rst,matrix_A[7012],matrix_B[12],mul_res1[7012]);
multi_7x28 multi_7x28_mod_7013(clk,rst,matrix_A[7013],matrix_B[13],mul_res1[7013]);
multi_7x28 multi_7x28_mod_7014(clk,rst,matrix_A[7014],matrix_B[14],mul_res1[7014]);
multi_7x28 multi_7x28_mod_7015(clk,rst,matrix_A[7015],matrix_B[15],mul_res1[7015]);
multi_7x28 multi_7x28_mod_7016(clk,rst,matrix_A[7016],matrix_B[16],mul_res1[7016]);
multi_7x28 multi_7x28_mod_7017(clk,rst,matrix_A[7017],matrix_B[17],mul_res1[7017]);
multi_7x28 multi_7x28_mod_7018(clk,rst,matrix_A[7018],matrix_B[18],mul_res1[7018]);
multi_7x28 multi_7x28_mod_7019(clk,rst,matrix_A[7019],matrix_B[19],mul_res1[7019]);
multi_7x28 multi_7x28_mod_7020(clk,rst,matrix_A[7020],matrix_B[20],mul_res1[7020]);
multi_7x28 multi_7x28_mod_7021(clk,rst,matrix_A[7021],matrix_B[21],mul_res1[7021]);
multi_7x28 multi_7x28_mod_7022(clk,rst,matrix_A[7022],matrix_B[22],mul_res1[7022]);
multi_7x28 multi_7x28_mod_7023(clk,rst,matrix_A[7023],matrix_B[23],mul_res1[7023]);
multi_7x28 multi_7x28_mod_7024(clk,rst,matrix_A[7024],matrix_B[24],mul_res1[7024]);
multi_7x28 multi_7x28_mod_7025(clk,rst,matrix_A[7025],matrix_B[25],mul_res1[7025]);
multi_7x28 multi_7x28_mod_7026(clk,rst,matrix_A[7026],matrix_B[26],mul_res1[7026]);
multi_7x28 multi_7x28_mod_7027(clk,rst,matrix_A[7027],matrix_B[27],mul_res1[7027]);
multi_7x28 multi_7x28_mod_7028(clk,rst,matrix_A[7028],matrix_B[28],mul_res1[7028]);
multi_7x28 multi_7x28_mod_7029(clk,rst,matrix_A[7029],matrix_B[29],mul_res1[7029]);
multi_7x28 multi_7x28_mod_7030(clk,rst,matrix_A[7030],matrix_B[30],mul_res1[7030]);
multi_7x28 multi_7x28_mod_7031(clk,rst,matrix_A[7031],matrix_B[31],mul_res1[7031]);
multi_7x28 multi_7x28_mod_7032(clk,rst,matrix_A[7032],matrix_B[32],mul_res1[7032]);
multi_7x28 multi_7x28_mod_7033(clk,rst,matrix_A[7033],matrix_B[33],mul_res1[7033]);
multi_7x28 multi_7x28_mod_7034(clk,rst,matrix_A[7034],matrix_B[34],mul_res1[7034]);
multi_7x28 multi_7x28_mod_7035(clk,rst,matrix_A[7035],matrix_B[35],mul_res1[7035]);
multi_7x28 multi_7x28_mod_7036(clk,rst,matrix_A[7036],matrix_B[36],mul_res1[7036]);
multi_7x28 multi_7x28_mod_7037(clk,rst,matrix_A[7037],matrix_B[37],mul_res1[7037]);
multi_7x28 multi_7x28_mod_7038(clk,rst,matrix_A[7038],matrix_B[38],mul_res1[7038]);
multi_7x28 multi_7x28_mod_7039(clk,rst,matrix_A[7039],matrix_B[39],mul_res1[7039]);
multi_7x28 multi_7x28_mod_7040(clk,rst,matrix_A[7040],matrix_B[40],mul_res1[7040]);
multi_7x28 multi_7x28_mod_7041(clk,rst,matrix_A[7041],matrix_B[41],mul_res1[7041]);
multi_7x28 multi_7x28_mod_7042(clk,rst,matrix_A[7042],matrix_B[42],mul_res1[7042]);
multi_7x28 multi_7x28_mod_7043(clk,rst,matrix_A[7043],matrix_B[43],mul_res1[7043]);
multi_7x28 multi_7x28_mod_7044(clk,rst,matrix_A[7044],matrix_B[44],mul_res1[7044]);
multi_7x28 multi_7x28_mod_7045(clk,rst,matrix_A[7045],matrix_B[45],mul_res1[7045]);
multi_7x28 multi_7x28_mod_7046(clk,rst,matrix_A[7046],matrix_B[46],mul_res1[7046]);
multi_7x28 multi_7x28_mod_7047(clk,rst,matrix_A[7047],matrix_B[47],mul_res1[7047]);
multi_7x28 multi_7x28_mod_7048(clk,rst,matrix_A[7048],matrix_B[48],mul_res1[7048]);
multi_7x28 multi_7x28_mod_7049(clk,rst,matrix_A[7049],matrix_B[49],mul_res1[7049]);
multi_7x28 multi_7x28_mod_7050(clk,rst,matrix_A[7050],matrix_B[50],mul_res1[7050]);
multi_7x28 multi_7x28_mod_7051(clk,rst,matrix_A[7051],matrix_B[51],mul_res1[7051]);
multi_7x28 multi_7x28_mod_7052(clk,rst,matrix_A[7052],matrix_B[52],mul_res1[7052]);
multi_7x28 multi_7x28_mod_7053(clk,rst,matrix_A[7053],matrix_B[53],mul_res1[7053]);
multi_7x28 multi_7x28_mod_7054(clk,rst,matrix_A[7054],matrix_B[54],mul_res1[7054]);
multi_7x28 multi_7x28_mod_7055(clk,rst,matrix_A[7055],matrix_B[55],mul_res1[7055]);
multi_7x28 multi_7x28_mod_7056(clk,rst,matrix_A[7056],matrix_B[56],mul_res1[7056]);
multi_7x28 multi_7x28_mod_7057(clk,rst,matrix_A[7057],matrix_B[57],mul_res1[7057]);
multi_7x28 multi_7x28_mod_7058(clk,rst,matrix_A[7058],matrix_B[58],mul_res1[7058]);
multi_7x28 multi_7x28_mod_7059(clk,rst,matrix_A[7059],matrix_B[59],mul_res1[7059]);
multi_7x28 multi_7x28_mod_7060(clk,rst,matrix_A[7060],matrix_B[60],mul_res1[7060]);
multi_7x28 multi_7x28_mod_7061(clk,rst,matrix_A[7061],matrix_B[61],mul_res1[7061]);
multi_7x28 multi_7x28_mod_7062(clk,rst,matrix_A[7062],matrix_B[62],mul_res1[7062]);
multi_7x28 multi_7x28_mod_7063(clk,rst,matrix_A[7063],matrix_B[63],mul_res1[7063]);
multi_7x28 multi_7x28_mod_7064(clk,rst,matrix_A[7064],matrix_B[64],mul_res1[7064]);
multi_7x28 multi_7x28_mod_7065(clk,rst,matrix_A[7065],matrix_B[65],mul_res1[7065]);
multi_7x28 multi_7x28_mod_7066(clk,rst,matrix_A[7066],matrix_B[66],mul_res1[7066]);
multi_7x28 multi_7x28_mod_7067(clk,rst,matrix_A[7067],matrix_B[67],mul_res1[7067]);
multi_7x28 multi_7x28_mod_7068(clk,rst,matrix_A[7068],matrix_B[68],mul_res1[7068]);
multi_7x28 multi_7x28_mod_7069(clk,rst,matrix_A[7069],matrix_B[69],mul_res1[7069]);
multi_7x28 multi_7x28_mod_7070(clk,rst,matrix_A[7070],matrix_B[70],mul_res1[7070]);
multi_7x28 multi_7x28_mod_7071(clk,rst,matrix_A[7071],matrix_B[71],mul_res1[7071]);
multi_7x28 multi_7x28_mod_7072(clk,rst,matrix_A[7072],matrix_B[72],mul_res1[7072]);
multi_7x28 multi_7x28_mod_7073(clk,rst,matrix_A[7073],matrix_B[73],mul_res1[7073]);
multi_7x28 multi_7x28_mod_7074(clk,rst,matrix_A[7074],matrix_B[74],mul_res1[7074]);
multi_7x28 multi_7x28_mod_7075(clk,rst,matrix_A[7075],matrix_B[75],mul_res1[7075]);
multi_7x28 multi_7x28_mod_7076(clk,rst,matrix_A[7076],matrix_B[76],mul_res1[7076]);
multi_7x28 multi_7x28_mod_7077(clk,rst,matrix_A[7077],matrix_B[77],mul_res1[7077]);
multi_7x28 multi_7x28_mod_7078(clk,rst,matrix_A[7078],matrix_B[78],mul_res1[7078]);
multi_7x28 multi_7x28_mod_7079(clk,rst,matrix_A[7079],matrix_B[79],mul_res1[7079]);
multi_7x28 multi_7x28_mod_7080(clk,rst,matrix_A[7080],matrix_B[80],mul_res1[7080]);
multi_7x28 multi_7x28_mod_7081(clk,rst,matrix_A[7081],matrix_B[81],mul_res1[7081]);
multi_7x28 multi_7x28_mod_7082(clk,rst,matrix_A[7082],matrix_B[82],mul_res1[7082]);
multi_7x28 multi_7x28_mod_7083(clk,rst,matrix_A[7083],matrix_B[83],mul_res1[7083]);
multi_7x28 multi_7x28_mod_7084(clk,rst,matrix_A[7084],matrix_B[84],mul_res1[7084]);
multi_7x28 multi_7x28_mod_7085(clk,rst,matrix_A[7085],matrix_B[85],mul_res1[7085]);
multi_7x28 multi_7x28_mod_7086(clk,rst,matrix_A[7086],matrix_B[86],mul_res1[7086]);
multi_7x28 multi_7x28_mod_7087(clk,rst,matrix_A[7087],matrix_B[87],mul_res1[7087]);
multi_7x28 multi_7x28_mod_7088(clk,rst,matrix_A[7088],matrix_B[88],mul_res1[7088]);
multi_7x28 multi_7x28_mod_7089(clk,rst,matrix_A[7089],matrix_B[89],mul_res1[7089]);
multi_7x28 multi_7x28_mod_7090(clk,rst,matrix_A[7090],matrix_B[90],mul_res1[7090]);
multi_7x28 multi_7x28_mod_7091(clk,rst,matrix_A[7091],matrix_B[91],mul_res1[7091]);
multi_7x28 multi_7x28_mod_7092(clk,rst,matrix_A[7092],matrix_B[92],mul_res1[7092]);
multi_7x28 multi_7x28_mod_7093(clk,rst,matrix_A[7093],matrix_B[93],mul_res1[7093]);
multi_7x28 multi_7x28_mod_7094(clk,rst,matrix_A[7094],matrix_B[94],mul_res1[7094]);
multi_7x28 multi_7x28_mod_7095(clk,rst,matrix_A[7095],matrix_B[95],mul_res1[7095]);
multi_7x28 multi_7x28_mod_7096(clk,rst,matrix_A[7096],matrix_B[96],mul_res1[7096]);
multi_7x28 multi_7x28_mod_7097(clk,rst,matrix_A[7097],matrix_B[97],mul_res1[7097]);
multi_7x28 multi_7x28_mod_7098(clk,rst,matrix_A[7098],matrix_B[98],mul_res1[7098]);
multi_7x28 multi_7x28_mod_7099(clk,rst,matrix_A[7099],matrix_B[99],mul_res1[7099]);
multi_7x28 multi_7x28_mod_7100(clk,rst,matrix_A[7100],matrix_B[100],mul_res1[7100]);
multi_7x28 multi_7x28_mod_7101(clk,rst,matrix_A[7101],matrix_B[101],mul_res1[7101]);
multi_7x28 multi_7x28_mod_7102(clk,rst,matrix_A[7102],matrix_B[102],mul_res1[7102]);
multi_7x28 multi_7x28_mod_7103(clk,rst,matrix_A[7103],matrix_B[103],mul_res1[7103]);
multi_7x28 multi_7x28_mod_7104(clk,rst,matrix_A[7104],matrix_B[104],mul_res1[7104]);
multi_7x28 multi_7x28_mod_7105(clk,rst,matrix_A[7105],matrix_B[105],mul_res1[7105]);
multi_7x28 multi_7x28_mod_7106(clk,rst,matrix_A[7106],matrix_B[106],mul_res1[7106]);
multi_7x28 multi_7x28_mod_7107(clk,rst,matrix_A[7107],matrix_B[107],mul_res1[7107]);
multi_7x28 multi_7x28_mod_7108(clk,rst,matrix_A[7108],matrix_B[108],mul_res1[7108]);
multi_7x28 multi_7x28_mod_7109(clk,rst,matrix_A[7109],matrix_B[109],mul_res1[7109]);
multi_7x28 multi_7x28_mod_7110(clk,rst,matrix_A[7110],matrix_B[110],mul_res1[7110]);
multi_7x28 multi_7x28_mod_7111(clk,rst,matrix_A[7111],matrix_B[111],mul_res1[7111]);
multi_7x28 multi_7x28_mod_7112(clk,rst,matrix_A[7112],matrix_B[112],mul_res1[7112]);
multi_7x28 multi_7x28_mod_7113(clk,rst,matrix_A[7113],matrix_B[113],mul_res1[7113]);
multi_7x28 multi_7x28_mod_7114(clk,rst,matrix_A[7114],matrix_B[114],mul_res1[7114]);
multi_7x28 multi_7x28_mod_7115(clk,rst,matrix_A[7115],matrix_B[115],mul_res1[7115]);
multi_7x28 multi_7x28_mod_7116(clk,rst,matrix_A[7116],matrix_B[116],mul_res1[7116]);
multi_7x28 multi_7x28_mod_7117(clk,rst,matrix_A[7117],matrix_B[117],mul_res1[7117]);
multi_7x28 multi_7x28_mod_7118(clk,rst,matrix_A[7118],matrix_B[118],mul_res1[7118]);
multi_7x28 multi_7x28_mod_7119(clk,rst,matrix_A[7119],matrix_B[119],mul_res1[7119]);
multi_7x28 multi_7x28_mod_7120(clk,rst,matrix_A[7120],matrix_B[120],mul_res1[7120]);
multi_7x28 multi_7x28_mod_7121(clk,rst,matrix_A[7121],matrix_B[121],mul_res1[7121]);
multi_7x28 multi_7x28_mod_7122(clk,rst,matrix_A[7122],matrix_B[122],mul_res1[7122]);
multi_7x28 multi_7x28_mod_7123(clk,rst,matrix_A[7123],matrix_B[123],mul_res1[7123]);
multi_7x28 multi_7x28_mod_7124(clk,rst,matrix_A[7124],matrix_B[124],mul_res1[7124]);
multi_7x28 multi_7x28_mod_7125(clk,rst,matrix_A[7125],matrix_B[125],mul_res1[7125]);
multi_7x28 multi_7x28_mod_7126(clk,rst,matrix_A[7126],matrix_B[126],mul_res1[7126]);
multi_7x28 multi_7x28_mod_7127(clk,rst,matrix_A[7127],matrix_B[127],mul_res1[7127]);
multi_7x28 multi_7x28_mod_7128(clk,rst,matrix_A[7128],matrix_B[128],mul_res1[7128]);
multi_7x28 multi_7x28_mod_7129(clk,rst,matrix_A[7129],matrix_B[129],mul_res1[7129]);
multi_7x28 multi_7x28_mod_7130(clk,rst,matrix_A[7130],matrix_B[130],mul_res1[7130]);
multi_7x28 multi_7x28_mod_7131(clk,rst,matrix_A[7131],matrix_B[131],mul_res1[7131]);
multi_7x28 multi_7x28_mod_7132(clk,rst,matrix_A[7132],matrix_B[132],mul_res1[7132]);
multi_7x28 multi_7x28_mod_7133(clk,rst,matrix_A[7133],matrix_B[133],mul_res1[7133]);
multi_7x28 multi_7x28_mod_7134(clk,rst,matrix_A[7134],matrix_B[134],mul_res1[7134]);
multi_7x28 multi_7x28_mod_7135(clk,rst,matrix_A[7135],matrix_B[135],mul_res1[7135]);
multi_7x28 multi_7x28_mod_7136(clk,rst,matrix_A[7136],matrix_B[136],mul_res1[7136]);
multi_7x28 multi_7x28_mod_7137(clk,rst,matrix_A[7137],matrix_B[137],mul_res1[7137]);
multi_7x28 multi_7x28_mod_7138(clk,rst,matrix_A[7138],matrix_B[138],mul_res1[7138]);
multi_7x28 multi_7x28_mod_7139(clk,rst,matrix_A[7139],matrix_B[139],mul_res1[7139]);
multi_7x28 multi_7x28_mod_7140(clk,rst,matrix_A[7140],matrix_B[140],mul_res1[7140]);
multi_7x28 multi_7x28_mod_7141(clk,rst,matrix_A[7141],matrix_B[141],mul_res1[7141]);
multi_7x28 multi_7x28_mod_7142(clk,rst,matrix_A[7142],matrix_B[142],mul_res1[7142]);
multi_7x28 multi_7x28_mod_7143(clk,rst,matrix_A[7143],matrix_B[143],mul_res1[7143]);
multi_7x28 multi_7x28_mod_7144(clk,rst,matrix_A[7144],matrix_B[144],mul_res1[7144]);
multi_7x28 multi_7x28_mod_7145(clk,rst,matrix_A[7145],matrix_B[145],mul_res1[7145]);
multi_7x28 multi_7x28_mod_7146(clk,rst,matrix_A[7146],matrix_B[146],mul_res1[7146]);
multi_7x28 multi_7x28_mod_7147(clk,rst,matrix_A[7147],matrix_B[147],mul_res1[7147]);
multi_7x28 multi_7x28_mod_7148(clk,rst,matrix_A[7148],matrix_B[148],mul_res1[7148]);
multi_7x28 multi_7x28_mod_7149(clk,rst,matrix_A[7149],matrix_B[149],mul_res1[7149]);
multi_7x28 multi_7x28_mod_7150(clk,rst,matrix_A[7150],matrix_B[150],mul_res1[7150]);
multi_7x28 multi_7x28_mod_7151(clk,rst,matrix_A[7151],matrix_B[151],mul_res1[7151]);
multi_7x28 multi_7x28_mod_7152(clk,rst,matrix_A[7152],matrix_B[152],mul_res1[7152]);
multi_7x28 multi_7x28_mod_7153(clk,rst,matrix_A[7153],matrix_B[153],mul_res1[7153]);
multi_7x28 multi_7x28_mod_7154(clk,rst,matrix_A[7154],matrix_B[154],mul_res1[7154]);
multi_7x28 multi_7x28_mod_7155(clk,rst,matrix_A[7155],matrix_B[155],mul_res1[7155]);
multi_7x28 multi_7x28_mod_7156(clk,rst,matrix_A[7156],matrix_B[156],mul_res1[7156]);
multi_7x28 multi_7x28_mod_7157(clk,rst,matrix_A[7157],matrix_B[157],mul_res1[7157]);
multi_7x28 multi_7x28_mod_7158(clk,rst,matrix_A[7158],matrix_B[158],mul_res1[7158]);
multi_7x28 multi_7x28_mod_7159(clk,rst,matrix_A[7159],matrix_B[159],mul_res1[7159]);
multi_7x28 multi_7x28_mod_7160(clk,rst,matrix_A[7160],matrix_B[160],mul_res1[7160]);
multi_7x28 multi_7x28_mod_7161(clk,rst,matrix_A[7161],matrix_B[161],mul_res1[7161]);
multi_7x28 multi_7x28_mod_7162(clk,rst,matrix_A[7162],matrix_B[162],mul_res1[7162]);
multi_7x28 multi_7x28_mod_7163(clk,rst,matrix_A[7163],matrix_B[163],mul_res1[7163]);
multi_7x28 multi_7x28_mod_7164(clk,rst,matrix_A[7164],matrix_B[164],mul_res1[7164]);
multi_7x28 multi_7x28_mod_7165(clk,rst,matrix_A[7165],matrix_B[165],mul_res1[7165]);
multi_7x28 multi_7x28_mod_7166(clk,rst,matrix_A[7166],matrix_B[166],mul_res1[7166]);
multi_7x28 multi_7x28_mod_7167(clk,rst,matrix_A[7167],matrix_B[167],mul_res1[7167]);
multi_7x28 multi_7x28_mod_7168(clk,rst,matrix_A[7168],matrix_B[168],mul_res1[7168]);
multi_7x28 multi_7x28_mod_7169(clk,rst,matrix_A[7169],matrix_B[169],mul_res1[7169]);
multi_7x28 multi_7x28_mod_7170(clk,rst,matrix_A[7170],matrix_B[170],mul_res1[7170]);
multi_7x28 multi_7x28_mod_7171(clk,rst,matrix_A[7171],matrix_B[171],mul_res1[7171]);
multi_7x28 multi_7x28_mod_7172(clk,rst,matrix_A[7172],matrix_B[172],mul_res1[7172]);
multi_7x28 multi_7x28_mod_7173(clk,rst,matrix_A[7173],matrix_B[173],mul_res1[7173]);
multi_7x28 multi_7x28_mod_7174(clk,rst,matrix_A[7174],matrix_B[174],mul_res1[7174]);
multi_7x28 multi_7x28_mod_7175(clk,rst,matrix_A[7175],matrix_B[175],mul_res1[7175]);
multi_7x28 multi_7x28_mod_7176(clk,rst,matrix_A[7176],matrix_B[176],mul_res1[7176]);
multi_7x28 multi_7x28_mod_7177(clk,rst,matrix_A[7177],matrix_B[177],mul_res1[7177]);
multi_7x28 multi_7x28_mod_7178(clk,rst,matrix_A[7178],matrix_B[178],mul_res1[7178]);
multi_7x28 multi_7x28_mod_7179(clk,rst,matrix_A[7179],matrix_B[179],mul_res1[7179]);
multi_7x28 multi_7x28_mod_7180(clk,rst,matrix_A[7180],matrix_B[180],mul_res1[7180]);
multi_7x28 multi_7x28_mod_7181(clk,rst,matrix_A[7181],matrix_B[181],mul_res1[7181]);
multi_7x28 multi_7x28_mod_7182(clk,rst,matrix_A[7182],matrix_B[182],mul_res1[7182]);
multi_7x28 multi_7x28_mod_7183(clk,rst,matrix_A[7183],matrix_B[183],mul_res1[7183]);
multi_7x28 multi_7x28_mod_7184(clk,rst,matrix_A[7184],matrix_B[184],mul_res1[7184]);
multi_7x28 multi_7x28_mod_7185(clk,rst,matrix_A[7185],matrix_B[185],mul_res1[7185]);
multi_7x28 multi_7x28_mod_7186(clk,rst,matrix_A[7186],matrix_B[186],mul_res1[7186]);
multi_7x28 multi_7x28_mod_7187(clk,rst,matrix_A[7187],matrix_B[187],mul_res1[7187]);
multi_7x28 multi_7x28_mod_7188(clk,rst,matrix_A[7188],matrix_B[188],mul_res1[7188]);
multi_7x28 multi_7x28_mod_7189(clk,rst,matrix_A[7189],matrix_B[189],mul_res1[7189]);
multi_7x28 multi_7x28_mod_7190(clk,rst,matrix_A[7190],matrix_B[190],mul_res1[7190]);
multi_7x28 multi_7x28_mod_7191(clk,rst,matrix_A[7191],matrix_B[191],mul_res1[7191]);
multi_7x28 multi_7x28_mod_7192(clk,rst,matrix_A[7192],matrix_B[192],mul_res1[7192]);
multi_7x28 multi_7x28_mod_7193(clk,rst,matrix_A[7193],matrix_B[193],mul_res1[7193]);
multi_7x28 multi_7x28_mod_7194(clk,rst,matrix_A[7194],matrix_B[194],mul_res1[7194]);
multi_7x28 multi_7x28_mod_7195(clk,rst,matrix_A[7195],matrix_B[195],mul_res1[7195]);
multi_7x28 multi_7x28_mod_7196(clk,rst,matrix_A[7196],matrix_B[196],mul_res1[7196]);
multi_7x28 multi_7x28_mod_7197(clk,rst,matrix_A[7197],matrix_B[197],mul_res1[7197]);
multi_7x28 multi_7x28_mod_7198(clk,rst,matrix_A[7198],matrix_B[198],mul_res1[7198]);
multi_7x28 multi_7x28_mod_7199(clk,rst,matrix_A[7199],matrix_B[199],mul_res1[7199]);
multi_7x28 multi_7x28_mod_7200(clk,rst,matrix_A[7200],matrix_B[0],mul_res1[7200]);
multi_7x28 multi_7x28_mod_7201(clk,rst,matrix_A[7201],matrix_B[1],mul_res1[7201]);
multi_7x28 multi_7x28_mod_7202(clk,rst,matrix_A[7202],matrix_B[2],mul_res1[7202]);
multi_7x28 multi_7x28_mod_7203(clk,rst,matrix_A[7203],matrix_B[3],mul_res1[7203]);
multi_7x28 multi_7x28_mod_7204(clk,rst,matrix_A[7204],matrix_B[4],mul_res1[7204]);
multi_7x28 multi_7x28_mod_7205(clk,rst,matrix_A[7205],matrix_B[5],mul_res1[7205]);
multi_7x28 multi_7x28_mod_7206(clk,rst,matrix_A[7206],matrix_B[6],mul_res1[7206]);
multi_7x28 multi_7x28_mod_7207(clk,rst,matrix_A[7207],matrix_B[7],mul_res1[7207]);
multi_7x28 multi_7x28_mod_7208(clk,rst,matrix_A[7208],matrix_B[8],mul_res1[7208]);
multi_7x28 multi_7x28_mod_7209(clk,rst,matrix_A[7209],matrix_B[9],mul_res1[7209]);
multi_7x28 multi_7x28_mod_7210(clk,rst,matrix_A[7210],matrix_B[10],mul_res1[7210]);
multi_7x28 multi_7x28_mod_7211(clk,rst,matrix_A[7211],matrix_B[11],mul_res1[7211]);
multi_7x28 multi_7x28_mod_7212(clk,rst,matrix_A[7212],matrix_B[12],mul_res1[7212]);
multi_7x28 multi_7x28_mod_7213(clk,rst,matrix_A[7213],matrix_B[13],mul_res1[7213]);
multi_7x28 multi_7x28_mod_7214(clk,rst,matrix_A[7214],matrix_B[14],mul_res1[7214]);
multi_7x28 multi_7x28_mod_7215(clk,rst,matrix_A[7215],matrix_B[15],mul_res1[7215]);
multi_7x28 multi_7x28_mod_7216(clk,rst,matrix_A[7216],matrix_B[16],mul_res1[7216]);
multi_7x28 multi_7x28_mod_7217(clk,rst,matrix_A[7217],matrix_B[17],mul_res1[7217]);
multi_7x28 multi_7x28_mod_7218(clk,rst,matrix_A[7218],matrix_B[18],mul_res1[7218]);
multi_7x28 multi_7x28_mod_7219(clk,rst,matrix_A[7219],matrix_B[19],mul_res1[7219]);
multi_7x28 multi_7x28_mod_7220(clk,rst,matrix_A[7220],matrix_B[20],mul_res1[7220]);
multi_7x28 multi_7x28_mod_7221(clk,rst,matrix_A[7221],matrix_B[21],mul_res1[7221]);
multi_7x28 multi_7x28_mod_7222(clk,rst,matrix_A[7222],matrix_B[22],mul_res1[7222]);
multi_7x28 multi_7x28_mod_7223(clk,rst,matrix_A[7223],matrix_B[23],mul_res1[7223]);
multi_7x28 multi_7x28_mod_7224(clk,rst,matrix_A[7224],matrix_B[24],mul_res1[7224]);
multi_7x28 multi_7x28_mod_7225(clk,rst,matrix_A[7225],matrix_B[25],mul_res1[7225]);
multi_7x28 multi_7x28_mod_7226(clk,rst,matrix_A[7226],matrix_B[26],mul_res1[7226]);
multi_7x28 multi_7x28_mod_7227(clk,rst,matrix_A[7227],matrix_B[27],mul_res1[7227]);
multi_7x28 multi_7x28_mod_7228(clk,rst,matrix_A[7228],matrix_B[28],mul_res1[7228]);
multi_7x28 multi_7x28_mod_7229(clk,rst,matrix_A[7229],matrix_B[29],mul_res1[7229]);
multi_7x28 multi_7x28_mod_7230(clk,rst,matrix_A[7230],matrix_B[30],mul_res1[7230]);
multi_7x28 multi_7x28_mod_7231(clk,rst,matrix_A[7231],matrix_B[31],mul_res1[7231]);
multi_7x28 multi_7x28_mod_7232(clk,rst,matrix_A[7232],matrix_B[32],mul_res1[7232]);
multi_7x28 multi_7x28_mod_7233(clk,rst,matrix_A[7233],matrix_B[33],mul_res1[7233]);
multi_7x28 multi_7x28_mod_7234(clk,rst,matrix_A[7234],matrix_B[34],mul_res1[7234]);
multi_7x28 multi_7x28_mod_7235(clk,rst,matrix_A[7235],matrix_B[35],mul_res1[7235]);
multi_7x28 multi_7x28_mod_7236(clk,rst,matrix_A[7236],matrix_B[36],mul_res1[7236]);
multi_7x28 multi_7x28_mod_7237(clk,rst,matrix_A[7237],matrix_B[37],mul_res1[7237]);
multi_7x28 multi_7x28_mod_7238(clk,rst,matrix_A[7238],matrix_B[38],mul_res1[7238]);
multi_7x28 multi_7x28_mod_7239(clk,rst,matrix_A[7239],matrix_B[39],mul_res1[7239]);
multi_7x28 multi_7x28_mod_7240(clk,rst,matrix_A[7240],matrix_B[40],mul_res1[7240]);
multi_7x28 multi_7x28_mod_7241(clk,rst,matrix_A[7241],matrix_B[41],mul_res1[7241]);
multi_7x28 multi_7x28_mod_7242(clk,rst,matrix_A[7242],matrix_B[42],mul_res1[7242]);
multi_7x28 multi_7x28_mod_7243(clk,rst,matrix_A[7243],matrix_B[43],mul_res1[7243]);
multi_7x28 multi_7x28_mod_7244(clk,rst,matrix_A[7244],matrix_B[44],mul_res1[7244]);
multi_7x28 multi_7x28_mod_7245(clk,rst,matrix_A[7245],matrix_B[45],mul_res1[7245]);
multi_7x28 multi_7x28_mod_7246(clk,rst,matrix_A[7246],matrix_B[46],mul_res1[7246]);
multi_7x28 multi_7x28_mod_7247(clk,rst,matrix_A[7247],matrix_B[47],mul_res1[7247]);
multi_7x28 multi_7x28_mod_7248(clk,rst,matrix_A[7248],matrix_B[48],mul_res1[7248]);
multi_7x28 multi_7x28_mod_7249(clk,rst,matrix_A[7249],matrix_B[49],mul_res1[7249]);
multi_7x28 multi_7x28_mod_7250(clk,rst,matrix_A[7250],matrix_B[50],mul_res1[7250]);
multi_7x28 multi_7x28_mod_7251(clk,rst,matrix_A[7251],matrix_B[51],mul_res1[7251]);
multi_7x28 multi_7x28_mod_7252(clk,rst,matrix_A[7252],matrix_B[52],mul_res1[7252]);
multi_7x28 multi_7x28_mod_7253(clk,rst,matrix_A[7253],matrix_B[53],mul_res1[7253]);
multi_7x28 multi_7x28_mod_7254(clk,rst,matrix_A[7254],matrix_B[54],mul_res1[7254]);
multi_7x28 multi_7x28_mod_7255(clk,rst,matrix_A[7255],matrix_B[55],mul_res1[7255]);
multi_7x28 multi_7x28_mod_7256(clk,rst,matrix_A[7256],matrix_B[56],mul_res1[7256]);
multi_7x28 multi_7x28_mod_7257(clk,rst,matrix_A[7257],matrix_B[57],mul_res1[7257]);
multi_7x28 multi_7x28_mod_7258(clk,rst,matrix_A[7258],matrix_B[58],mul_res1[7258]);
multi_7x28 multi_7x28_mod_7259(clk,rst,matrix_A[7259],matrix_B[59],mul_res1[7259]);
multi_7x28 multi_7x28_mod_7260(clk,rst,matrix_A[7260],matrix_B[60],mul_res1[7260]);
multi_7x28 multi_7x28_mod_7261(clk,rst,matrix_A[7261],matrix_B[61],mul_res1[7261]);
multi_7x28 multi_7x28_mod_7262(clk,rst,matrix_A[7262],matrix_B[62],mul_res1[7262]);
multi_7x28 multi_7x28_mod_7263(clk,rst,matrix_A[7263],matrix_B[63],mul_res1[7263]);
multi_7x28 multi_7x28_mod_7264(clk,rst,matrix_A[7264],matrix_B[64],mul_res1[7264]);
multi_7x28 multi_7x28_mod_7265(clk,rst,matrix_A[7265],matrix_B[65],mul_res1[7265]);
multi_7x28 multi_7x28_mod_7266(clk,rst,matrix_A[7266],matrix_B[66],mul_res1[7266]);
multi_7x28 multi_7x28_mod_7267(clk,rst,matrix_A[7267],matrix_B[67],mul_res1[7267]);
multi_7x28 multi_7x28_mod_7268(clk,rst,matrix_A[7268],matrix_B[68],mul_res1[7268]);
multi_7x28 multi_7x28_mod_7269(clk,rst,matrix_A[7269],matrix_B[69],mul_res1[7269]);
multi_7x28 multi_7x28_mod_7270(clk,rst,matrix_A[7270],matrix_B[70],mul_res1[7270]);
multi_7x28 multi_7x28_mod_7271(clk,rst,matrix_A[7271],matrix_B[71],mul_res1[7271]);
multi_7x28 multi_7x28_mod_7272(clk,rst,matrix_A[7272],matrix_B[72],mul_res1[7272]);
multi_7x28 multi_7x28_mod_7273(clk,rst,matrix_A[7273],matrix_B[73],mul_res1[7273]);
multi_7x28 multi_7x28_mod_7274(clk,rst,matrix_A[7274],matrix_B[74],mul_res1[7274]);
multi_7x28 multi_7x28_mod_7275(clk,rst,matrix_A[7275],matrix_B[75],mul_res1[7275]);
multi_7x28 multi_7x28_mod_7276(clk,rst,matrix_A[7276],matrix_B[76],mul_res1[7276]);
multi_7x28 multi_7x28_mod_7277(clk,rst,matrix_A[7277],matrix_B[77],mul_res1[7277]);
multi_7x28 multi_7x28_mod_7278(clk,rst,matrix_A[7278],matrix_B[78],mul_res1[7278]);
multi_7x28 multi_7x28_mod_7279(clk,rst,matrix_A[7279],matrix_B[79],mul_res1[7279]);
multi_7x28 multi_7x28_mod_7280(clk,rst,matrix_A[7280],matrix_B[80],mul_res1[7280]);
multi_7x28 multi_7x28_mod_7281(clk,rst,matrix_A[7281],matrix_B[81],mul_res1[7281]);
multi_7x28 multi_7x28_mod_7282(clk,rst,matrix_A[7282],matrix_B[82],mul_res1[7282]);
multi_7x28 multi_7x28_mod_7283(clk,rst,matrix_A[7283],matrix_B[83],mul_res1[7283]);
multi_7x28 multi_7x28_mod_7284(clk,rst,matrix_A[7284],matrix_B[84],mul_res1[7284]);
multi_7x28 multi_7x28_mod_7285(clk,rst,matrix_A[7285],matrix_B[85],mul_res1[7285]);
multi_7x28 multi_7x28_mod_7286(clk,rst,matrix_A[7286],matrix_B[86],mul_res1[7286]);
multi_7x28 multi_7x28_mod_7287(clk,rst,matrix_A[7287],matrix_B[87],mul_res1[7287]);
multi_7x28 multi_7x28_mod_7288(clk,rst,matrix_A[7288],matrix_B[88],mul_res1[7288]);
multi_7x28 multi_7x28_mod_7289(clk,rst,matrix_A[7289],matrix_B[89],mul_res1[7289]);
multi_7x28 multi_7x28_mod_7290(clk,rst,matrix_A[7290],matrix_B[90],mul_res1[7290]);
multi_7x28 multi_7x28_mod_7291(clk,rst,matrix_A[7291],matrix_B[91],mul_res1[7291]);
multi_7x28 multi_7x28_mod_7292(clk,rst,matrix_A[7292],matrix_B[92],mul_res1[7292]);
multi_7x28 multi_7x28_mod_7293(clk,rst,matrix_A[7293],matrix_B[93],mul_res1[7293]);
multi_7x28 multi_7x28_mod_7294(clk,rst,matrix_A[7294],matrix_B[94],mul_res1[7294]);
multi_7x28 multi_7x28_mod_7295(clk,rst,matrix_A[7295],matrix_B[95],mul_res1[7295]);
multi_7x28 multi_7x28_mod_7296(clk,rst,matrix_A[7296],matrix_B[96],mul_res1[7296]);
multi_7x28 multi_7x28_mod_7297(clk,rst,matrix_A[7297],matrix_B[97],mul_res1[7297]);
multi_7x28 multi_7x28_mod_7298(clk,rst,matrix_A[7298],matrix_B[98],mul_res1[7298]);
multi_7x28 multi_7x28_mod_7299(clk,rst,matrix_A[7299],matrix_B[99],mul_res1[7299]);
multi_7x28 multi_7x28_mod_7300(clk,rst,matrix_A[7300],matrix_B[100],mul_res1[7300]);
multi_7x28 multi_7x28_mod_7301(clk,rst,matrix_A[7301],matrix_B[101],mul_res1[7301]);
multi_7x28 multi_7x28_mod_7302(clk,rst,matrix_A[7302],matrix_B[102],mul_res1[7302]);
multi_7x28 multi_7x28_mod_7303(clk,rst,matrix_A[7303],matrix_B[103],mul_res1[7303]);
multi_7x28 multi_7x28_mod_7304(clk,rst,matrix_A[7304],matrix_B[104],mul_res1[7304]);
multi_7x28 multi_7x28_mod_7305(clk,rst,matrix_A[7305],matrix_B[105],mul_res1[7305]);
multi_7x28 multi_7x28_mod_7306(clk,rst,matrix_A[7306],matrix_B[106],mul_res1[7306]);
multi_7x28 multi_7x28_mod_7307(clk,rst,matrix_A[7307],matrix_B[107],mul_res1[7307]);
multi_7x28 multi_7x28_mod_7308(clk,rst,matrix_A[7308],matrix_B[108],mul_res1[7308]);
multi_7x28 multi_7x28_mod_7309(clk,rst,matrix_A[7309],matrix_B[109],mul_res1[7309]);
multi_7x28 multi_7x28_mod_7310(clk,rst,matrix_A[7310],matrix_B[110],mul_res1[7310]);
multi_7x28 multi_7x28_mod_7311(clk,rst,matrix_A[7311],matrix_B[111],mul_res1[7311]);
multi_7x28 multi_7x28_mod_7312(clk,rst,matrix_A[7312],matrix_B[112],mul_res1[7312]);
multi_7x28 multi_7x28_mod_7313(clk,rst,matrix_A[7313],matrix_B[113],mul_res1[7313]);
multi_7x28 multi_7x28_mod_7314(clk,rst,matrix_A[7314],matrix_B[114],mul_res1[7314]);
multi_7x28 multi_7x28_mod_7315(clk,rst,matrix_A[7315],matrix_B[115],mul_res1[7315]);
multi_7x28 multi_7x28_mod_7316(clk,rst,matrix_A[7316],matrix_B[116],mul_res1[7316]);
multi_7x28 multi_7x28_mod_7317(clk,rst,matrix_A[7317],matrix_B[117],mul_res1[7317]);
multi_7x28 multi_7x28_mod_7318(clk,rst,matrix_A[7318],matrix_B[118],mul_res1[7318]);
multi_7x28 multi_7x28_mod_7319(clk,rst,matrix_A[7319],matrix_B[119],mul_res1[7319]);
multi_7x28 multi_7x28_mod_7320(clk,rst,matrix_A[7320],matrix_B[120],mul_res1[7320]);
multi_7x28 multi_7x28_mod_7321(clk,rst,matrix_A[7321],matrix_B[121],mul_res1[7321]);
multi_7x28 multi_7x28_mod_7322(clk,rst,matrix_A[7322],matrix_B[122],mul_res1[7322]);
multi_7x28 multi_7x28_mod_7323(clk,rst,matrix_A[7323],matrix_B[123],mul_res1[7323]);
multi_7x28 multi_7x28_mod_7324(clk,rst,matrix_A[7324],matrix_B[124],mul_res1[7324]);
multi_7x28 multi_7x28_mod_7325(clk,rst,matrix_A[7325],matrix_B[125],mul_res1[7325]);
multi_7x28 multi_7x28_mod_7326(clk,rst,matrix_A[7326],matrix_B[126],mul_res1[7326]);
multi_7x28 multi_7x28_mod_7327(clk,rst,matrix_A[7327],matrix_B[127],mul_res1[7327]);
multi_7x28 multi_7x28_mod_7328(clk,rst,matrix_A[7328],matrix_B[128],mul_res1[7328]);
multi_7x28 multi_7x28_mod_7329(clk,rst,matrix_A[7329],matrix_B[129],mul_res1[7329]);
multi_7x28 multi_7x28_mod_7330(clk,rst,matrix_A[7330],matrix_B[130],mul_res1[7330]);
multi_7x28 multi_7x28_mod_7331(clk,rst,matrix_A[7331],matrix_B[131],mul_res1[7331]);
multi_7x28 multi_7x28_mod_7332(clk,rst,matrix_A[7332],matrix_B[132],mul_res1[7332]);
multi_7x28 multi_7x28_mod_7333(clk,rst,matrix_A[7333],matrix_B[133],mul_res1[7333]);
multi_7x28 multi_7x28_mod_7334(clk,rst,matrix_A[7334],matrix_B[134],mul_res1[7334]);
multi_7x28 multi_7x28_mod_7335(clk,rst,matrix_A[7335],matrix_B[135],mul_res1[7335]);
multi_7x28 multi_7x28_mod_7336(clk,rst,matrix_A[7336],matrix_B[136],mul_res1[7336]);
multi_7x28 multi_7x28_mod_7337(clk,rst,matrix_A[7337],matrix_B[137],mul_res1[7337]);
multi_7x28 multi_7x28_mod_7338(clk,rst,matrix_A[7338],matrix_B[138],mul_res1[7338]);
multi_7x28 multi_7x28_mod_7339(clk,rst,matrix_A[7339],matrix_B[139],mul_res1[7339]);
multi_7x28 multi_7x28_mod_7340(clk,rst,matrix_A[7340],matrix_B[140],mul_res1[7340]);
multi_7x28 multi_7x28_mod_7341(clk,rst,matrix_A[7341],matrix_B[141],mul_res1[7341]);
multi_7x28 multi_7x28_mod_7342(clk,rst,matrix_A[7342],matrix_B[142],mul_res1[7342]);
multi_7x28 multi_7x28_mod_7343(clk,rst,matrix_A[7343],matrix_B[143],mul_res1[7343]);
multi_7x28 multi_7x28_mod_7344(clk,rst,matrix_A[7344],matrix_B[144],mul_res1[7344]);
multi_7x28 multi_7x28_mod_7345(clk,rst,matrix_A[7345],matrix_B[145],mul_res1[7345]);
multi_7x28 multi_7x28_mod_7346(clk,rst,matrix_A[7346],matrix_B[146],mul_res1[7346]);
multi_7x28 multi_7x28_mod_7347(clk,rst,matrix_A[7347],matrix_B[147],mul_res1[7347]);
multi_7x28 multi_7x28_mod_7348(clk,rst,matrix_A[7348],matrix_B[148],mul_res1[7348]);
multi_7x28 multi_7x28_mod_7349(clk,rst,matrix_A[7349],matrix_B[149],mul_res1[7349]);
multi_7x28 multi_7x28_mod_7350(clk,rst,matrix_A[7350],matrix_B[150],mul_res1[7350]);
multi_7x28 multi_7x28_mod_7351(clk,rst,matrix_A[7351],matrix_B[151],mul_res1[7351]);
multi_7x28 multi_7x28_mod_7352(clk,rst,matrix_A[7352],matrix_B[152],mul_res1[7352]);
multi_7x28 multi_7x28_mod_7353(clk,rst,matrix_A[7353],matrix_B[153],mul_res1[7353]);
multi_7x28 multi_7x28_mod_7354(clk,rst,matrix_A[7354],matrix_B[154],mul_res1[7354]);
multi_7x28 multi_7x28_mod_7355(clk,rst,matrix_A[7355],matrix_B[155],mul_res1[7355]);
multi_7x28 multi_7x28_mod_7356(clk,rst,matrix_A[7356],matrix_B[156],mul_res1[7356]);
multi_7x28 multi_7x28_mod_7357(clk,rst,matrix_A[7357],matrix_B[157],mul_res1[7357]);
multi_7x28 multi_7x28_mod_7358(clk,rst,matrix_A[7358],matrix_B[158],mul_res1[7358]);
multi_7x28 multi_7x28_mod_7359(clk,rst,matrix_A[7359],matrix_B[159],mul_res1[7359]);
multi_7x28 multi_7x28_mod_7360(clk,rst,matrix_A[7360],matrix_B[160],mul_res1[7360]);
multi_7x28 multi_7x28_mod_7361(clk,rst,matrix_A[7361],matrix_B[161],mul_res1[7361]);
multi_7x28 multi_7x28_mod_7362(clk,rst,matrix_A[7362],matrix_B[162],mul_res1[7362]);
multi_7x28 multi_7x28_mod_7363(clk,rst,matrix_A[7363],matrix_B[163],mul_res1[7363]);
multi_7x28 multi_7x28_mod_7364(clk,rst,matrix_A[7364],matrix_B[164],mul_res1[7364]);
multi_7x28 multi_7x28_mod_7365(clk,rst,matrix_A[7365],matrix_B[165],mul_res1[7365]);
multi_7x28 multi_7x28_mod_7366(clk,rst,matrix_A[7366],matrix_B[166],mul_res1[7366]);
multi_7x28 multi_7x28_mod_7367(clk,rst,matrix_A[7367],matrix_B[167],mul_res1[7367]);
multi_7x28 multi_7x28_mod_7368(clk,rst,matrix_A[7368],matrix_B[168],mul_res1[7368]);
multi_7x28 multi_7x28_mod_7369(clk,rst,matrix_A[7369],matrix_B[169],mul_res1[7369]);
multi_7x28 multi_7x28_mod_7370(clk,rst,matrix_A[7370],matrix_B[170],mul_res1[7370]);
multi_7x28 multi_7x28_mod_7371(clk,rst,matrix_A[7371],matrix_B[171],mul_res1[7371]);
multi_7x28 multi_7x28_mod_7372(clk,rst,matrix_A[7372],matrix_B[172],mul_res1[7372]);
multi_7x28 multi_7x28_mod_7373(clk,rst,matrix_A[7373],matrix_B[173],mul_res1[7373]);
multi_7x28 multi_7x28_mod_7374(clk,rst,matrix_A[7374],matrix_B[174],mul_res1[7374]);
multi_7x28 multi_7x28_mod_7375(clk,rst,matrix_A[7375],matrix_B[175],mul_res1[7375]);
multi_7x28 multi_7x28_mod_7376(clk,rst,matrix_A[7376],matrix_B[176],mul_res1[7376]);
multi_7x28 multi_7x28_mod_7377(clk,rst,matrix_A[7377],matrix_B[177],mul_res1[7377]);
multi_7x28 multi_7x28_mod_7378(clk,rst,matrix_A[7378],matrix_B[178],mul_res1[7378]);
multi_7x28 multi_7x28_mod_7379(clk,rst,matrix_A[7379],matrix_B[179],mul_res1[7379]);
multi_7x28 multi_7x28_mod_7380(clk,rst,matrix_A[7380],matrix_B[180],mul_res1[7380]);
multi_7x28 multi_7x28_mod_7381(clk,rst,matrix_A[7381],matrix_B[181],mul_res1[7381]);
multi_7x28 multi_7x28_mod_7382(clk,rst,matrix_A[7382],matrix_B[182],mul_res1[7382]);
multi_7x28 multi_7x28_mod_7383(clk,rst,matrix_A[7383],matrix_B[183],mul_res1[7383]);
multi_7x28 multi_7x28_mod_7384(clk,rst,matrix_A[7384],matrix_B[184],mul_res1[7384]);
multi_7x28 multi_7x28_mod_7385(clk,rst,matrix_A[7385],matrix_B[185],mul_res1[7385]);
multi_7x28 multi_7x28_mod_7386(clk,rst,matrix_A[7386],matrix_B[186],mul_res1[7386]);
multi_7x28 multi_7x28_mod_7387(clk,rst,matrix_A[7387],matrix_B[187],mul_res1[7387]);
multi_7x28 multi_7x28_mod_7388(clk,rst,matrix_A[7388],matrix_B[188],mul_res1[7388]);
multi_7x28 multi_7x28_mod_7389(clk,rst,matrix_A[7389],matrix_B[189],mul_res1[7389]);
multi_7x28 multi_7x28_mod_7390(clk,rst,matrix_A[7390],matrix_B[190],mul_res1[7390]);
multi_7x28 multi_7x28_mod_7391(clk,rst,matrix_A[7391],matrix_B[191],mul_res1[7391]);
multi_7x28 multi_7x28_mod_7392(clk,rst,matrix_A[7392],matrix_B[192],mul_res1[7392]);
multi_7x28 multi_7x28_mod_7393(clk,rst,matrix_A[7393],matrix_B[193],mul_res1[7393]);
multi_7x28 multi_7x28_mod_7394(clk,rst,matrix_A[7394],matrix_B[194],mul_res1[7394]);
multi_7x28 multi_7x28_mod_7395(clk,rst,matrix_A[7395],matrix_B[195],mul_res1[7395]);
multi_7x28 multi_7x28_mod_7396(clk,rst,matrix_A[7396],matrix_B[196],mul_res1[7396]);
multi_7x28 multi_7x28_mod_7397(clk,rst,matrix_A[7397],matrix_B[197],mul_res1[7397]);
multi_7x28 multi_7x28_mod_7398(clk,rst,matrix_A[7398],matrix_B[198],mul_res1[7398]);
multi_7x28 multi_7x28_mod_7399(clk,rst,matrix_A[7399],matrix_B[199],mul_res1[7399]);
multi_7x28 multi_7x28_mod_7400(clk,rst,matrix_A[7400],matrix_B[0],mul_res1[7400]);
multi_7x28 multi_7x28_mod_7401(clk,rst,matrix_A[7401],matrix_B[1],mul_res1[7401]);
multi_7x28 multi_7x28_mod_7402(clk,rst,matrix_A[7402],matrix_B[2],mul_res1[7402]);
multi_7x28 multi_7x28_mod_7403(clk,rst,matrix_A[7403],matrix_B[3],mul_res1[7403]);
multi_7x28 multi_7x28_mod_7404(clk,rst,matrix_A[7404],matrix_B[4],mul_res1[7404]);
multi_7x28 multi_7x28_mod_7405(clk,rst,matrix_A[7405],matrix_B[5],mul_res1[7405]);
multi_7x28 multi_7x28_mod_7406(clk,rst,matrix_A[7406],matrix_B[6],mul_res1[7406]);
multi_7x28 multi_7x28_mod_7407(clk,rst,matrix_A[7407],matrix_B[7],mul_res1[7407]);
multi_7x28 multi_7x28_mod_7408(clk,rst,matrix_A[7408],matrix_B[8],mul_res1[7408]);
multi_7x28 multi_7x28_mod_7409(clk,rst,matrix_A[7409],matrix_B[9],mul_res1[7409]);
multi_7x28 multi_7x28_mod_7410(clk,rst,matrix_A[7410],matrix_B[10],mul_res1[7410]);
multi_7x28 multi_7x28_mod_7411(clk,rst,matrix_A[7411],matrix_B[11],mul_res1[7411]);
multi_7x28 multi_7x28_mod_7412(clk,rst,matrix_A[7412],matrix_B[12],mul_res1[7412]);
multi_7x28 multi_7x28_mod_7413(clk,rst,matrix_A[7413],matrix_B[13],mul_res1[7413]);
multi_7x28 multi_7x28_mod_7414(clk,rst,matrix_A[7414],matrix_B[14],mul_res1[7414]);
multi_7x28 multi_7x28_mod_7415(clk,rst,matrix_A[7415],matrix_B[15],mul_res1[7415]);
multi_7x28 multi_7x28_mod_7416(clk,rst,matrix_A[7416],matrix_B[16],mul_res1[7416]);
multi_7x28 multi_7x28_mod_7417(clk,rst,matrix_A[7417],matrix_B[17],mul_res1[7417]);
multi_7x28 multi_7x28_mod_7418(clk,rst,matrix_A[7418],matrix_B[18],mul_res1[7418]);
multi_7x28 multi_7x28_mod_7419(clk,rst,matrix_A[7419],matrix_B[19],mul_res1[7419]);
multi_7x28 multi_7x28_mod_7420(clk,rst,matrix_A[7420],matrix_B[20],mul_res1[7420]);
multi_7x28 multi_7x28_mod_7421(clk,rst,matrix_A[7421],matrix_B[21],mul_res1[7421]);
multi_7x28 multi_7x28_mod_7422(clk,rst,matrix_A[7422],matrix_B[22],mul_res1[7422]);
multi_7x28 multi_7x28_mod_7423(clk,rst,matrix_A[7423],matrix_B[23],mul_res1[7423]);
multi_7x28 multi_7x28_mod_7424(clk,rst,matrix_A[7424],matrix_B[24],mul_res1[7424]);
multi_7x28 multi_7x28_mod_7425(clk,rst,matrix_A[7425],matrix_B[25],mul_res1[7425]);
multi_7x28 multi_7x28_mod_7426(clk,rst,matrix_A[7426],matrix_B[26],mul_res1[7426]);
multi_7x28 multi_7x28_mod_7427(clk,rst,matrix_A[7427],matrix_B[27],mul_res1[7427]);
multi_7x28 multi_7x28_mod_7428(clk,rst,matrix_A[7428],matrix_B[28],mul_res1[7428]);
multi_7x28 multi_7x28_mod_7429(clk,rst,matrix_A[7429],matrix_B[29],mul_res1[7429]);
multi_7x28 multi_7x28_mod_7430(clk,rst,matrix_A[7430],matrix_B[30],mul_res1[7430]);
multi_7x28 multi_7x28_mod_7431(clk,rst,matrix_A[7431],matrix_B[31],mul_res1[7431]);
multi_7x28 multi_7x28_mod_7432(clk,rst,matrix_A[7432],matrix_B[32],mul_res1[7432]);
multi_7x28 multi_7x28_mod_7433(clk,rst,matrix_A[7433],matrix_B[33],mul_res1[7433]);
multi_7x28 multi_7x28_mod_7434(clk,rst,matrix_A[7434],matrix_B[34],mul_res1[7434]);
multi_7x28 multi_7x28_mod_7435(clk,rst,matrix_A[7435],matrix_B[35],mul_res1[7435]);
multi_7x28 multi_7x28_mod_7436(clk,rst,matrix_A[7436],matrix_B[36],mul_res1[7436]);
multi_7x28 multi_7x28_mod_7437(clk,rst,matrix_A[7437],matrix_B[37],mul_res1[7437]);
multi_7x28 multi_7x28_mod_7438(clk,rst,matrix_A[7438],matrix_B[38],mul_res1[7438]);
multi_7x28 multi_7x28_mod_7439(clk,rst,matrix_A[7439],matrix_B[39],mul_res1[7439]);
multi_7x28 multi_7x28_mod_7440(clk,rst,matrix_A[7440],matrix_B[40],mul_res1[7440]);
multi_7x28 multi_7x28_mod_7441(clk,rst,matrix_A[7441],matrix_B[41],mul_res1[7441]);
multi_7x28 multi_7x28_mod_7442(clk,rst,matrix_A[7442],matrix_B[42],mul_res1[7442]);
multi_7x28 multi_7x28_mod_7443(clk,rst,matrix_A[7443],matrix_B[43],mul_res1[7443]);
multi_7x28 multi_7x28_mod_7444(clk,rst,matrix_A[7444],matrix_B[44],mul_res1[7444]);
multi_7x28 multi_7x28_mod_7445(clk,rst,matrix_A[7445],matrix_B[45],mul_res1[7445]);
multi_7x28 multi_7x28_mod_7446(clk,rst,matrix_A[7446],matrix_B[46],mul_res1[7446]);
multi_7x28 multi_7x28_mod_7447(clk,rst,matrix_A[7447],matrix_B[47],mul_res1[7447]);
multi_7x28 multi_7x28_mod_7448(clk,rst,matrix_A[7448],matrix_B[48],mul_res1[7448]);
multi_7x28 multi_7x28_mod_7449(clk,rst,matrix_A[7449],matrix_B[49],mul_res1[7449]);
multi_7x28 multi_7x28_mod_7450(clk,rst,matrix_A[7450],matrix_B[50],mul_res1[7450]);
multi_7x28 multi_7x28_mod_7451(clk,rst,matrix_A[7451],matrix_B[51],mul_res1[7451]);
multi_7x28 multi_7x28_mod_7452(clk,rst,matrix_A[7452],matrix_B[52],mul_res1[7452]);
multi_7x28 multi_7x28_mod_7453(clk,rst,matrix_A[7453],matrix_B[53],mul_res1[7453]);
multi_7x28 multi_7x28_mod_7454(clk,rst,matrix_A[7454],matrix_B[54],mul_res1[7454]);
multi_7x28 multi_7x28_mod_7455(clk,rst,matrix_A[7455],matrix_B[55],mul_res1[7455]);
multi_7x28 multi_7x28_mod_7456(clk,rst,matrix_A[7456],matrix_B[56],mul_res1[7456]);
multi_7x28 multi_7x28_mod_7457(clk,rst,matrix_A[7457],matrix_B[57],mul_res1[7457]);
multi_7x28 multi_7x28_mod_7458(clk,rst,matrix_A[7458],matrix_B[58],mul_res1[7458]);
multi_7x28 multi_7x28_mod_7459(clk,rst,matrix_A[7459],matrix_B[59],mul_res1[7459]);
multi_7x28 multi_7x28_mod_7460(clk,rst,matrix_A[7460],matrix_B[60],mul_res1[7460]);
multi_7x28 multi_7x28_mod_7461(clk,rst,matrix_A[7461],matrix_B[61],mul_res1[7461]);
multi_7x28 multi_7x28_mod_7462(clk,rst,matrix_A[7462],matrix_B[62],mul_res1[7462]);
multi_7x28 multi_7x28_mod_7463(clk,rst,matrix_A[7463],matrix_B[63],mul_res1[7463]);
multi_7x28 multi_7x28_mod_7464(clk,rst,matrix_A[7464],matrix_B[64],mul_res1[7464]);
multi_7x28 multi_7x28_mod_7465(clk,rst,matrix_A[7465],matrix_B[65],mul_res1[7465]);
multi_7x28 multi_7x28_mod_7466(clk,rst,matrix_A[7466],matrix_B[66],mul_res1[7466]);
multi_7x28 multi_7x28_mod_7467(clk,rst,matrix_A[7467],matrix_B[67],mul_res1[7467]);
multi_7x28 multi_7x28_mod_7468(clk,rst,matrix_A[7468],matrix_B[68],mul_res1[7468]);
multi_7x28 multi_7x28_mod_7469(clk,rst,matrix_A[7469],matrix_B[69],mul_res1[7469]);
multi_7x28 multi_7x28_mod_7470(clk,rst,matrix_A[7470],matrix_B[70],mul_res1[7470]);
multi_7x28 multi_7x28_mod_7471(clk,rst,matrix_A[7471],matrix_B[71],mul_res1[7471]);
multi_7x28 multi_7x28_mod_7472(clk,rst,matrix_A[7472],matrix_B[72],mul_res1[7472]);
multi_7x28 multi_7x28_mod_7473(clk,rst,matrix_A[7473],matrix_B[73],mul_res1[7473]);
multi_7x28 multi_7x28_mod_7474(clk,rst,matrix_A[7474],matrix_B[74],mul_res1[7474]);
multi_7x28 multi_7x28_mod_7475(clk,rst,matrix_A[7475],matrix_B[75],mul_res1[7475]);
multi_7x28 multi_7x28_mod_7476(clk,rst,matrix_A[7476],matrix_B[76],mul_res1[7476]);
multi_7x28 multi_7x28_mod_7477(clk,rst,matrix_A[7477],matrix_B[77],mul_res1[7477]);
multi_7x28 multi_7x28_mod_7478(clk,rst,matrix_A[7478],matrix_B[78],mul_res1[7478]);
multi_7x28 multi_7x28_mod_7479(clk,rst,matrix_A[7479],matrix_B[79],mul_res1[7479]);
multi_7x28 multi_7x28_mod_7480(clk,rst,matrix_A[7480],matrix_B[80],mul_res1[7480]);
multi_7x28 multi_7x28_mod_7481(clk,rst,matrix_A[7481],matrix_B[81],mul_res1[7481]);
multi_7x28 multi_7x28_mod_7482(clk,rst,matrix_A[7482],matrix_B[82],mul_res1[7482]);
multi_7x28 multi_7x28_mod_7483(clk,rst,matrix_A[7483],matrix_B[83],mul_res1[7483]);
multi_7x28 multi_7x28_mod_7484(clk,rst,matrix_A[7484],matrix_B[84],mul_res1[7484]);
multi_7x28 multi_7x28_mod_7485(clk,rst,matrix_A[7485],matrix_B[85],mul_res1[7485]);
multi_7x28 multi_7x28_mod_7486(clk,rst,matrix_A[7486],matrix_B[86],mul_res1[7486]);
multi_7x28 multi_7x28_mod_7487(clk,rst,matrix_A[7487],matrix_B[87],mul_res1[7487]);
multi_7x28 multi_7x28_mod_7488(clk,rst,matrix_A[7488],matrix_B[88],mul_res1[7488]);
multi_7x28 multi_7x28_mod_7489(clk,rst,matrix_A[7489],matrix_B[89],mul_res1[7489]);
multi_7x28 multi_7x28_mod_7490(clk,rst,matrix_A[7490],matrix_B[90],mul_res1[7490]);
multi_7x28 multi_7x28_mod_7491(clk,rst,matrix_A[7491],matrix_B[91],mul_res1[7491]);
multi_7x28 multi_7x28_mod_7492(clk,rst,matrix_A[7492],matrix_B[92],mul_res1[7492]);
multi_7x28 multi_7x28_mod_7493(clk,rst,matrix_A[7493],matrix_B[93],mul_res1[7493]);
multi_7x28 multi_7x28_mod_7494(clk,rst,matrix_A[7494],matrix_B[94],mul_res1[7494]);
multi_7x28 multi_7x28_mod_7495(clk,rst,matrix_A[7495],matrix_B[95],mul_res1[7495]);
multi_7x28 multi_7x28_mod_7496(clk,rst,matrix_A[7496],matrix_B[96],mul_res1[7496]);
multi_7x28 multi_7x28_mod_7497(clk,rst,matrix_A[7497],matrix_B[97],mul_res1[7497]);
multi_7x28 multi_7x28_mod_7498(clk,rst,matrix_A[7498],matrix_B[98],mul_res1[7498]);
multi_7x28 multi_7x28_mod_7499(clk,rst,matrix_A[7499],matrix_B[99],mul_res1[7499]);
multi_7x28 multi_7x28_mod_7500(clk,rst,matrix_A[7500],matrix_B[100],mul_res1[7500]);
multi_7x28 multi_7x28_mod_7501(clk,rst,matrix_A[7501],matrix_B[101],mul_res1[7501]);
multi_7x28 multi_7x28_mod_7502(clk,rst,matrix_A[7502],matrix_B[102],mul_res1[7502]);
multi_7x28 multi_7x28_mod_7503(clk,rst,matrix_A[7503],matrix_B[103],mul_res1[7503]);
multi_7x28 multi_7x28_mod_7504(clk,rst,matrix_A[7504],matrix_B[104],mul_res1[7504]);
multi_7x28 multi_7x28_mod_7505(clk,rst,matrix_A[7505],matrix_B[105],mul_res1[7505]);
multi_7x28 multi_7x28_mod_7506(clk,rst,matrix_A[7506],matrix_B[106],mul_res1[7506]);
multi_7x28 multi_7x28_mod_7507(clk,rst,matrix_A[7507],matrix_B[107],mul_res1[7507]);
multi_7x28 multi_7x28_mod_7508(clk,rst,matrix_A[7508],matrix_B[108],mul_res1[7508]);
multi_7x28 multi_7x28_mod_7509(clk,rst,matrix_A[7509],matrix_B[109],mul_res1[7509]);
multi_7x28 multi_7x28_mod_7510(clk,rst,matrix_A[7510],matrix_B[110],mul_res1[7510]);
multi_7x28 multi_7x28_mod_7511(clk,rst,matrix_A[7511],matrix_B[111],mul_res1[7511]);
multi_7x28 multi_7x28_mod_7512(clk,rst,matrix_A[7512],matrix_B[112],mul_res1[7512]);
multi_7x28 multi_7x28_mod_7513(clk,rst,matrix_A[7513],matrix_B[113],mul_res1[7513]);
multi_7x28 multi_7x28_mod_7514(clk,rst,matrix_A[7514],matrix_B[114],mul_res1[7514]);
multi_7x28 multi_7x28_mod_7515(clk,rst,matrix_A[7515],matrix_B[115],mul_res1[7515]);
multi_7x28 multi_7x28_mod_7516(clk,rst,matrix_A[7516],matrix_B[116],mul_res1[7516]);
multi_7x28 multi_7x28_mod_7517(clk,rst,matrix_A[7517],matrix_B[117],mul_res1[7517]);
multi_7x28 multi_7x28_mod_7518(clk,rst,matrix_A[7518],matrix_B[118],mul_res1[7518]);
multi_7x28 multi_7x28_mod_7519(clk,rst,matrix_A[7519],matrix_B[119],mul_res1[7519]);
multi_7x28 multi_7x28_mod_7520(clk,rst,matrix_A[7520],matrix_B[120],mul_res1[7520]);
multi_7x28 multi_7x28_mod_7521(clk,rst,matrix_A[7521],matrix_B[121],mul_res1[7521]);
multi_7x28 multi_7x28_mod_7522(clk,rst,matrix_A[7522],matrix_B[122],mul_res1[7522]);
multi_7x28 multi_7x28_mod_7523(clk,rst,matrix_A[7523],matrix_B[123],mul_res1[7523]);
multi_7x28 multi_7x28_mod_7524(clk,rst,matrix_A[7524],matrix_B[124],mul_res1[7524]);
multi_7x28 multi_7x28_mod_7525(clk,rst,matrix_A[7525],matrix_B[125],mul_res1[7525]);
multi_7x28 multi_7x28_mod_7526(clk,rst,matrix_A[7526],matrix_B[126],mul_res1[7526]);
multi_7x28 multi_7x28_mod_7527(clk,rst,matrix_A[7527],matrix_B[127],mul_res1[7527]);
multi_7x28 multi_7x28_mod_7528(clk,rst,matrix_A[7528],matrix_B[128],mul_res1[7528]);
multi_7x28 multi_7x28_mod_7529(clk,rst,matrix_A[7529],matrix_B[129],mul_res1[7529]);
multi_7x28 multi_7x28_mod_7530(clk,rst,matrix_A[7530],matrix_B[130],mul_res1[7530]);
multi_7x28 multi_7x28_mod_7531(clk,rst,matrix_A[7531],matrix_B[131],mul_res1[7531]);
multi_7x28 multi_7x28_mod_7532(clk,rst,matrix_A[7532],matrix_B[132],mul_res1[7532]);
multi_7x28 multi_7x28_mod_7533(clk,rst,matrix_A[7533],matrix_B[133],mul_res1[7533]);
multi_7x28 multi_7x28_mod_7534(clk,rst,matrix_A[7534],matrix_B[134],mul_res1[7534]);
multi_7x28 multi_7x28_mod_7535(clk,rst,matrix_A[7535],matrix_B[135],mul_res1[7535]);
multi_7x28 multi_7x28_mod_7536(clk,rst,matrix_A[7536],matrix_B[136],mul_res1[7536]);
multi_7x28 multi_7x28_mod_7537(clk,rst,matrix_A[7537],matrix_B[137],mul_res1[7537]);
multi_7x28 multi_7x28_mod_7538(clk,rst,matrix_A[7538],matrix_B[138],mul_res1[7538]);
multi_7x28 multi_7x28_mod_7539(clk,rst,matrix_A[7539],matrix_B[139],mul_res1[7539]);
multi_7x28 multi_7x28_mod_7540(clk,rst,matrix_A[7540],matrix_B[140],mul_res1[7540]);
multi_7x28 multi_7x28_mod_7541(clk,rst,matrix_A[7541],matrix_B[141],mul_res1[7541]);
multi_7x28 multi_7x28_mod_7542(clk,rst,matrix_A[7542],matrix_B[142],mul_res1[7542]);
multi_7x28 multi_7x28_mod_7543(clk,rst,matrix_A[7543],matrix_B[143],mul_res1[7543]);
multi_7x28 multi_7x28_mod_7544(clk,rst,matrix_A[7544],matrix_B[144],mul_res1[7544]);
multi_7x28 multi_7x28_mod_7545(clk,rst,matrix_A[7545],matrix_B[145],mul_res1[7545]);
multi_7x28 multi_7x28_mod_7546(clk,rst,matrix_A[7546],matrix_B[146],mul_res1[7546]);
multi_7x28 multi_7x28_mod_7547(clk,rst,matrix_A[7547],matrix_B[147],mul_res1[7547]);
multi_7x28 multi_7x28_mod_7548(clk,rst,matrix_A[7548],matrix_B[148],mul_res1[7548]);
multi_7x28 multi_7x28_mod_7549(clk,rst,matrix_A[7549],matrix_B[149],mul_res1[7549]);
multi_7x28 multi_7x28_mod_7550(clk,rst,matrix_A[7550],matrix_B[150],mul_res1[7550]);
multi_7x28 multi_7x28_mod_7551(clk,rst,matrix_A[7551],matrix_B[151],mul_res1[7551]);
multi_7x28 multi_7x28_mod_7552(clk,rst,matrix_A[7552],matrix_B[152],mul_res1[7552]);
multi_7x28 multi_7x28_mod_7553(clk,rst,matrix_A[7553],matrix_B[153],mul_res1[7553]);
multi_7x28 multi_7x28_mod_7554(clk,rst,matrix_A[7554],matrix_B[154],mul_res1[7554]);
multi_7x28 multi_7x28_mod_7555(clk,rst,matrix_A[7555],matrix_B[155],mul_res1[7555]);
multi_7x28 multi_7x28_mod_7556(clk,rst,matrix_A[7556],matrix_B[156],mul_res1[7556]);
multi_7x28 multi_7x28_mod_7557(clk,rst,matrix_A[7557],matrix_B[157],mul_res1[7557]);
multi_7x28 multi_7x28_mod_7558(clk,rst,matrix_A[7558],matrix_B[158],mul_res1[7558]);
multi_7x28 multi_7x28_mod_7559(clk,rst,matrix_A[7559],matrix_B[159],mul_res1[7559]);
multi_7x28 multi_7x28_mod_7560(clk,rst,matrix_A[7560],matrix_B[160],mul_res1[7560]);
multi_7x28 multi_7x28_mod_7561(clk,rst,matrix_A[7561],matrix_B[161],mul_res1[7561]);
multi_7x28 multi_7x28_mod_7562(clk,rst,matrix_A[7562],matrix_B[162],mul_res1[7562]);
multi_7x28 multi_7x28_mod_7563(clk,rst,matrix_A[7563],matrix_B[163],mul_res1[7563]);
multi_7x28 multi_7x28_mod_7564(clk,rst,matrix_A[7564],matrix_B[164],mul_res1[7564]);
multi_7x28 multi_7x28_mod_7565(clk,rst,matrix_A[7565],matrix_B[165],mul_res1[7565]);
multi_7x28 multi_7x28_mod_7566(clk,rst,matrix_A[7566],matrix_B[166],mul_res1[7566]);
multi_7x28 multi_7x28_mod_7567(clk,rst,matrix_A[7567],matrix_B[167],mul_res1[7567]);
multi_7x28 multi_7x28_mod_7568(clk,rst,matrix_A[7568],matrix_B[168],mul_res1[7568]);
multi_7x28 multi_7x28_mod_7569(clk,rst,matrix_A[7569],matrix_B[169],mul_res1[7569]);
multi_7x28 multi_7x28_mod_7570(clk,rst,matrix_A[7570],matrix_B[170],mul_res1[7570]);
multi_7x28 multi_7x28_mod_7571(clk,rst,matrix_A[7571],matrix_B[171],mul_res1[7571]);
multi_7x28 multi_7x28_mod_7572(clk,rst,matrix_A[7572],matrix_B[172],mul_res1[7572]);
multi_7x28 multi_7x28_mod_7573(clk,rst,matrix_A[7573],matrix_B[173],mul_res1[7573]);
multi_7x28 multi_7x28_mod_7574(clk,rst,matrix_A[7574],matrix_B[174],mul_res1[7574]);
multi_7x28 multi_7x28_mod_7575(clk,rst,matrix_A[7575],matrix_B[175],mul_res1[7575]);
multi_7x28 multi_7x28_mod_7576(clk,rst,matrix_A[7576],matrix_B[176],mul_res1[7576]);
multi_7x28 multi_7x28_mod_7577(clk,rst,matrix_A[7577],matrix_B[177],mul_res1[7577]);
multi_7x28 multi_7x28_mod_7578(clk,rst,matrix_A[7578],matrix_B[178],mul_res1[7578]);
multi_7x28 multi_7x28_mod_7579(clk,rst,matrix_A[7579],matrix_B[179],mul_res1[7579]);
multi_7x28 multi_7x28_mod_7580(clk,rst,matrix_A[7580],matrix_B[180],mul_res1[7580]);
multi_7x28 multi_7x28_mod_7581(clk,rst,matrix_A[7581],matrix_B[181],mul_res1[7581]);
multi_7x28 multi_7x28_mod_7582(clk,rst,matrix_A[7582],matrix_B[182],mul_res1[7582]);
multi_7x28 multi_7x28_mod_7583(clk,rst,matrix_A[7583],matrix_B[183],mul_res1[7583]);
multi_7x28 multi_7x28_mod_7584(clk,rst,matrix_A[7584],matrix_B[184],mul_res1[7584]);
multi_7x28 multi_7x28_mod_7585(clk,rst,matrix_A[7585],matrix_B[185],mul_res1[7585]);
multi_7x28 multi_7x28_mod_7586(clk,rst,matrix_A[7586],matrix_B[186],mul_res1[7586]);
multi_7x28 multi_7x28_mod_7587(clk,rst,matrix_A[7587],matrix_B[187],mul_res1[7587]);
multi_7x28 multi_7x28_mod_7588(clk,rst,matrix_A[7588],matrix_B[188],mul_res1[7588]);
multi_7x28 multi_7x28_mod_7589(clk,rst,matrix_A[7589],matrix_B[189],mul_res1[7589]);
multi_7x28 multi_7x28_mod_7590(clk,rst,matrix_A[7590],matrix_B[190],mul_res1[7590]);
multi_7x28 multi_7x28_mod_7591(clk,rst,matrix_A[7591],matrix_B[191],mul_res1[7591]);
multi_7x28 multi_7x28_mod_7592(clk,rst,matrix_A[7592],matrix_B[192],mul_res1[7592]);
multi_7x28 multi_7x28_mod_7593(clk,rst,matrix_A[7593],matrix_B[193],mul_res1[7593]);
multi_7x28 multi_7x28_mod_7594(clk,rst,matrix_A[7594],matrix_B[194],mul_res1[7594]);
multi_7x28 multi_7x28_mod_7595(clk,rst,matrix_A[7595],matrix_B[195],mul_res1[7595]);
multi_7x28 multi_7x28_mod_7596(clk,rst,matrix_A[7596],matrix_B[196],mul_res1[7596]);
multi_7x28 multi_7x28_mod_7597(clk,rst,matrix_A[7597],matrix_B[197],mul_res1[7597]);
multi_7x28 multi_7x28_mod_7598(clk,rst,matrix_A[7598],matrix_B[198],mul_res1[7598]);
multi_7x28 multi_7x28_mod_7599(clk,rst,matrix_A[7599],matrix_B[199],mul_res1[7599]);
multi_7x28 multi_7x28_mod_7600(clk,rst,matrix_A[7600],matrix_B[0],mul_res1[7600]);
multi_7x28 multi_7x28_mod_7601(clk,rst,matrix_A[7601],matrix_B[1],mul_res1[7601]);
multi_7x28 multi_7x28_mod_7602(clk,rst,matrix_A[7602],matrix_B[2],mul_res1[7602]);
multi_7x28 multi_7x28_mod_7603(clk,rst,matrix_A[7603],matrix_B[3],mul_res1[7603]);
multi_7x28 multi_7x28_mod_7604(clk,rst,matrix_A[7604],matrix_B[4],mul_res1[7604]);
multi_7x28 multi_7x28_mod_7605(clk,rst,matrix_A[7605],matrix_B[5],mul_res1[7605]);
multi_7x28 multi_7x28_mod_7606(clk,rst,matrix_A[7606],matrix_B[6],mul_res1[7606]);
multi_7x28 multi_7x28_mod_7607(clk,rst,matrix_A[7607],matrix_B[7],mul_res1[7607]);
multi_7x28 multi_7x28_mod_7608(clk,rst,matrix_A[7608],matrix_B[8],mul_res1[7608]);
multi_7x28 multi_7x28_mod_7609(clk,rst,matrix_A[7609],matrix_B[9],mul_res1[7609]);
multi_7x28 multi_7x28_mod_7610(clk,rst,matrix_A[7610],matrix_B[10],mul_res1[7610]);
multi_7x28 multi_7x28_mod_7611(clk,rst,matrix_A[7611],matrix_B[11],mul_res1[7611]);
multi_7x28 multi_7x28_mod_7612(clk,rst,matrix_A[7612],matrix_B[12],mul_res1[7612]);
multi_7x28 multi_7x28_mod_7613(clk,rst,matrix_A[7613],matrix_B[13],mul_res1[7613]);
multi_7x28 multi_7x28_mod_7614(clk,rst,matrix_A[7614],matrix_B[14],mul_res1[7614]);
multi_7x28 multi_7x28_mod_7615(clk,rst,matrix_A[7615],matrix_B[15],mul_res1[7615]);
multi_7x28 multi_7x28_mod_7616(clk,rst,matrix_A[7616],matrix_B[16],mul_res1[7616]);
multi_7x28 multi_7x28_mod_7617(clk,rst,matrix_A[7617],matrix_B[17],mul_res1[7617]);
multi_7x28 multi_7x28_mod_7618(clk,rst,matrix_A[7618],matrix_B[18],mul_res1[7618]);
multi_7x28 multi_7x28_mod_7619(clk,rst,matrix_A[7619],matrix_B[19],mul_res1[7619]);
multi_7x28 multi_7x28_mod_7620(clk,rst,matrix_A[7620],matrix_B[20],mul_res1[7620]);
multi_7x28 multi_7x28_mod_7621(clk,rst,matrix_A[7621],matrix_B[21],mul_res1[7621]);
multi_7x28 multi_7x28_mod_7622(clk,rst,matrix_A[7622],matrix_B[22],mul_res1[7622]);
multi_7x28 multi_7x28_mod_7623(clk,rst,matrix_A[7623],matrix_B[23],mul_res1[7623]);
multi_7x28 multi_7x28_mod_7624(clk,rst,matrix_A[7624],matrix_B[24],mul_res1[7624]);
multi_7x28 multi_7x28_mod_7625(clk,rst,matrix_A[7625],matrix_B[25],mul_res1[7625]);
multi_7x28 multi_7x28_mod_7626(clk,rst,matrix_A[7626],matrix_B[26],mul_res1[7626]);
multi_7x28 multi_7x28_mod_7627(clk,rst,matrix_A[7627],matrix_B[27],mul_res1[7627]);
multi_7x28 multi_7x28_mod_7628(clk,rst,matrix_A[7628],matrix_B[28],mul_res1[7628]);
multi_7x28 multi_7x28_mod_7629(clk,rst,matrix_A[7629],matrix_B[29],mul_res1[7629]);
multi_7x28 multi_7x28_mod_7630(clk,rst,matrix_A[7630],matrix_B[30],mul_res1[7630]);
multi_7x28 multi_7x28_mod_7631(clk,rst,matrix_A[7631],matrix_B[31],mul_res1[7631]);
multi_7x28 multi_7x28_mod_7632(clk,rst,matrix_A[7632],matrix_B[32],mul_res1[7632]);
multi_7x28 multi_7x28_mod_7633(clk,rst,matrix_A[7633],matrix_B[33],mul_res1[7633]);
multi_7x28 multi_7x28_mod_7634(clk,rst,matrix_A[7634],matrix_B[34],mul_res1[7634]);
multi_7x28 multi_7x28_mod_7635(clk,rst,matrix_A[7635],matrix_B[35],mul_res1[7635]);
multi_7x28 multi_7x28_mod_7636(clk,rst,matrix_A[7636],matrix_B[36],mul_res1[7636]);
multi_7x28 multi_7x28_mod_7637(clk,rst,matrix_A[7637],matrix_B[37],mul_res1[7637]);
multi_7x28 multi_7x28_mod_7638(clk,rst,matrix_A[7638],matrix_B[38],mul_res1[7638]);
multi_7x28 multi_7x28_mod_7639(clk,rst,matrix_A[7639],matrix_B[39],mul_res1[7639]);
multi_7x28 multi_7x28_mod_7640(clk,rst,matrix_A[7640],matrix_B[40],mul_res1[7640]);
multi_7x28 multi_7x28_mod_7641(clk,rst,matrix_A[7641],matrix_B[41],mul_res1[7641]);
multi_7x28 multi_7x28_mod_7642(clk,rst,matrix_A[7642],matrix_B[42],mul_res1[7642]);
multi_7x28 multi_7x28_mod_7643(clk,rst,matrix_A[7643],matrix_B[43],mul_res1[7643]);
multi_7x28 multi_7x28_mod_7644(clk,rst,matrix_A[7644],matrix_B[44],mul_res1[7644]);
multi_7x28 multi_7x28_mod_7645(clk,rst,matrix_A[7645],matrix_B[45],mul_res1[7645]);
multi_7x28 multi_7x28_mod_7646(clk,rst,matrix_A[7646],matrix_B[46],mul_res1[7646]);
multi_7x28 multi_7x28_mod_7647(clk,rst,matrix_A[7647],matrix_B[47],mul_res1[7647]);
multi_7x28 multi_7x28_mod_7648(clk,rst,matrix_A[7648],matrix_B[48],mul_res1[7648]);
multi_7x28 multi_7x28_mod_7649(clk,rst,matrix_A[7649],matrix_B[49],mul_res1[7649]);
multi_7x28 multi_7x28_mod_7650(clk,rst,matrix_A[7650],matrix_B[50],mul_res1[7650]);
multi_7x28 multi_7x28_mod_7651(clk,rst,matrix_A[7651],matrix_B[51],mul_res1[7651]);
multi_7x28 multi_7x28_mod_7652(clk,rst,matrix_A[7652],matrix_B[52],mul_res1[7652]);
multi_7x28 multi_7x28_mod_7653(clk,rst,matrix_A[7653],matrix_B[53],mul_res1[7653]);
multi_7x28 multi_7x28_mod_7654(clk,rst,matrix_A[7654],matrix_B[54],mul_res1[7654]);
multi_7x28 multi_7x28_mod_7655(clk,rst,matrix_A[7655],matrix_B[55],mul_res1[7655]);
multi_7x28 multi_7x28_mod_7656(clk,rst,matrix_A[7656],matrix_B[56],mul_res1[7656]);
multi_7x28 multi_7x28_mod_7657(clk,rst,matrix_A[7657],matrix_B[57],mul_res1[7657]);
multi_7x28 multi_7x28_mod_7658(clk,rst,matrix_A[7658],matrix_B[58],mul_res1[7658]);
multi_7x28 multi_7x28_mod_7659(clk,rst,matrix_A[7659],matrix_B[59],mul_res1[7659]);
multi_7x28 multi_7x28_mod_7660(clk,rst,matrix_A[7660],matrix_B[60],mul_res1[7660]);
multi_7x28 multi_7x28_mod_7661(clk,rst,matrix_A[7661],matrix_B[61],mul_res1[7661]);
multi_7x28 multi_7x28_mod_7662(clk,rst,matrix_A[7662],matrix_B[62],mul_res1[7662]);
multi_7x28 multi_7x28_mod_7663(clk,rst,matrix_A[7663],matrix_B[63],mul_res1[7663]);
multi_7x28 multi_7x28_mod_7664(clk,rst,matrix_A[7664],matrix_B[64],mul_res1[7664]);
multi_7x28 multi_7x28_mod_7665(clk,rst,matrix_A[7665],matrix_B[65],mul_res1[7665]);
multi_7x28 multi_7x28_mod_7666(clk,rst,matrix_A[7666],matrix_B[66],mul_res1[7666]);
multi_7x28 multi_7x28_mod_7667(clk,rst,matrix_A[7667],matrix_B[67],mul_res1[7667]);
multi_7x28 multi_7x28_mod_7668(clk,rst,matrix_A[7668],matrix_B[68],mul_res1[7668]);
multi_7x28 multi_7x28_mod_7669(clk,rst,matrix_A[7669],matrix_B[69],mul_res1[7669]);
multi_7x28 multi_7x28_mod_7670(clk,rst,matrix_A[7670],matrix_B[70],mul_res1[7670]);
multi_7x28 multi_7x28_mod_7671(clk,rst,matrix_A[7671],matrix_B[71],mul_res1[7671]);
multi_7x28 multi_7x28_mod_7672(clk,rst,matrix_A[7672],matrix_B[72],mul_res1[7672]);
multi_7x28 multi_7x28_mod_7673(clk,rst,matrix_A[7673],matrix_B[73],mul_res1[7673]);
multi_7x28 multi_7x28_mod_7674(clk,rst,matrix_A[7674],matrix_B[74],mul_res1[7674]);
multi_7x28 multi_7x28_mod_7675(clk,rst,matrix_A[7675],matrix_B[75],mul_res1[7675]);
multi_7x28 multi_7x28_mod_7676(clk,rst,matrix_A[7676],matrix_B[76],mul_res1[7676]);
multi_7x28 multi_7x28_mod_7677(clk,rst,matrix_A[7677],matrix_B[77],mul_res1[7677]);
multi_7x28 multi_7x28_mod_7678(clk,rst,matrix_A[7678],matrix_B[78],mul_res1[7678]);
multi_7x28 multi_7x28_mod_7679(clk,rst,matrix_A[7679],matrix_B[79],mul_res1[7679]);
multi_7x28 multi_7x28_mod_7680(clk,rst,matrix_A[7680],matrix_B[80],mul_res1[7680]);
multi_7x28 multi_7x28_mod_7681(clk,rst,matrix_A[7681],matrix_B[81],mul_res1[7681]);
multi_7x28 multi_7x28_mod_7682(clk,rst,matrix_A[7682],matrix_B[82],mul_res1[7682]);
multi_7x28 multi_7x28_mod_7683(clk,rst,matrix_A[7683],matrix_B[83],mul_res1[7683]);
multi_7x28 multi_7x28_mod_7684(clk,rst,matrix_A[7684],matrix_B[84],mul_res1[7684]);
multi_7x28 multi_7x28_mod_7685(clk,rst,matrix_A[7685],matrix_B[85],mul_res1[7685]);
multi_7x28 multi_7x28_mod_7686(clk,rst,matrix_A[7686],matrix_B[86],mul_res1[7686]);
multi_7x28 multi_7x28_mod_7687(clk,rst,matrix_A[7687],matrix_B[87],mul_res1[7687]);
multi_7x28 multi_7x28_mod_7688(clk,rst,matrix_A[7688],matrix_B[88],mul_res1[7688]);
multi_7x28 multi_7x28_mod_7689(clk,rst,matrix_A[7689],matrix_B[89],mul_res1[7689]);
multi_7x28 multi_7x28_mod_7690(clk,rst,matrix_A[7690],matrix_B[90],mul_res1[7690]);
multi_7x28 multi_7x28_mod_7691(clk,rst,matrix_A[7691],matrix_B[91],mul_res1[7691]);
multi_7x28 multi_7x28_mod_7692(clk,rst,matrix_A[7692],matrix_B[92],mul_res1[7692]);
multi_7x28 multi_7x28_mod_7693(clk,rst,matrix_A[7693],matrix_B[93],mul_res1[7693]);
multi_7x28 multi_7x28_mod_7694(clk,rst,matrix_A[7694],matrix_B[94],mul_res1[7694]);
multi_7x28 multi_7x28_mod_7695(clk,rst,matrix_A[7695],matrix_B[95],mul_res1[7695]);
multi_7x28 multi_7x28_mod_7696(clk,rst,matrix_A[7696],matrix_B[96],mul_res1[7696]);
multi_7x28 multi_7x28_mod_7697(clk,rst,matrix_A[7697],matrix_B[97],mul_res1[7697]);
multi_7x28 multi_7x28_mod_7698(clk,rst,matrix_A[7698],matrix_B[98],mul_res1[7698]);
multi_7x28 multi_7x28_mod_7699(clk,rst,matrix_A[7699],matrix_B[99],mul_res1[7699]);
multi_7x28 multi_7x28_mod_7700(clk,rst,matrix_A[7700],matrix_B[100],mul_res1[7700]);
multi_7x28 multi_7x28_mod_7701(clk,rst,matrix_A[7701],matrix_B[101],mul_res1[7701]);
multi_7x28 multi_7x28_mod_7702(clk,rst,matrix_A[7702],matrix_B[102],mul_res1[7702]);
multi_7x28 multi_7x28_mod_7703(clk,rst,matrix_A[7703],matrix_B[103],mul_res1[7703]);
multi_7x28 multi_7x28_mod_7704(clk,rst,matrix_A[7704],matrix_B[104],mul_res1[7704]);
multi_7x28 multi_7x28_mod_7705(clk,rst,matrix_A[7705],matrix_B[105],mul_res1[7705]);
multi_7x28 multi_7x28_mod_7706(clk,rst,matrix_A[7706],matrix_B[106],mul_res1[7706]);
multi_7x28 multi_7x28_mod_7707(clk,rst,matrix_A[7707],matrix_B[107],mul_res1[7707]);
multi_7x28 multi_7x28_mod_7708(clk,rst,matrix_A[7708],matrix_B[108],mul_res1[7708]);
multi_7x28 multi_7x28_mod_7709(clk,rst,matrix_A[7709],matrix_B[109],mul_res1[7709]);
multi_7x28 multi_7x28_mod_7710(clk,rst,matrix_A[7710],matrix_B[110],mul_res1[7710]);
multi_7x28 multi_7x28_mod_7711(clk,rst,matrix_A[7711],matrix_B[111],mul_res1[7711]);
multi_7x28 multi_7x28_mod_7712(clk,rst,matrix_A[7712],matrix_B[112],mul_res1[7712]);
multi_7x28 multi_7x28_mod_7713(clk,rst,matrix_A[7713],matrix_B[113],mul_res1[7713]);
multi_7x28 multi_7x28_mod_7714(clk,rst,matrix_A[7714],matrix_B[114],mul_res1[7714]);
multi_7x28 multi_7x28_mod_7715(clk,rst,matrix_A[7715],matrix_B[115],mul_res1[7715]);
multi_7x28 multi_7x28_mod_7716(clk,rst,matrix_A[7716],matrix_B[116],mul_res1[7716]);
multi_7x28 multi_7x28_mod_7717(clk,rst,matrix_A[7717],matrix_B[117],mul_res1[7717]);
multi_7x28 multi_7x28_mod_7718(clk,rst,matrix_A[7718],matrix_B[118],mul_res1[7718]);
multi_7x28 multi_7x28_mod_7719(clk,rst,matrix_A[7719],matrix_B[119],mul_res1[7719]);
multi_7x28 multi_7x28_mod_7720(clk,rst,matrix_A[7720],matrix_B[120],mul_res1[7720]);
multi_7x28 multi_7x28_mod_7721(clk,rst,matrix_A[7721],matrix_B[121],mul_res1[7721]);
multi_7x28 multi_7x28_mod_7722(clk,rst,matrix_A[7722],matrix_B[122],mul_res1[7722]);
multi_7x28 multi_7x28_mod_7723(clk,rst,matrix_A[7723],matrix_B[123],mul_res1[7723]);
multi_7x28 multi_7x28_mod_7724(clk,rst,matrix_A[7724],matrix_B[124],mul_res1[7724]);
multi_7x28 multi_7x28_mod_7725(clk,rst,matrix_A[7725],matrix_B[125],mul_res1[7725]);
multi_7x28 multi_7x28_mod_7726(clk,rst,matrix_A[7726],matrix_B[126],mul_res1[7726]);
multi_7x28 multi_7x28_mod_7727(clk,rst,matrix_A[7727],matrix_B[127],mul_res1[7727]);
multi_7x28 multi_7x28_mod_7728(clk,rst,matrix_A[7728],matrix_B[128],mul_res1[7728]);
multi_7x28 multi_7x28_mod_7729(clk,rst,matrix_A[7729],matrix_B[129],mul_res1[7729]);
multi_7x28 multi_7x28_mod_7730(clk,rst,matrix_A[7730],matrix_B[130],mul_res1[7730]);
multi_7x28 multi_7x28_mod_7731(clk,rst,matrix_A[7731],matrix_B[131],mul_res1[7731]);
multi_7x28 multi_7x28_mod_7732(clk,rst,matrix_A[7732],matrix_B[132],mul_res1[7732]);
multi_7x28 multi_7x28_mod_7733(clk,rst,matrix_A[7733],matrix_B[133],mul_res1[7733]);
multi_7x28 multi_7x28_mod_7734(clk,rst,matrix_A[7734],matrix_B[134],mul_res1[7734]);
multi_7x28 multi_7x28_mod_7735(clk,rst,matrix_A[7735],matrix_B[135],mul_res1[7735]);
multi_7x28 multi_7x28_mod_7736(clk,rst,matrix_A[7736],matrix_B[136],mul_res1[7736]);
multi_7x28 multi_7x28_mod_7737(clk,rst,matrix_A[7737],matrix_B[137],mul_res1[7737]);
multi_7x28 multi_7x28_mod_7738(clk,rst,matrix_A[7738],matrix_B[138],mul_res1[7738]);
multi_7x28 multi_7x28_mod_7739(clk,rst,matrix_A[7739],matrix_B[139],mul_res1[7739]);
multi_7x28 multi_7x28_mod_7740(clk,rst,matrix_A[7740],matrix_B[140],mul_res1[7740]);
multi_7x28 multi_7x28_mod_7741(clk,rst,matrix_A[7741],matrix_B[141],mul_res1[7741]);
multi_7x28 multi_7x28_mod_7742(clk,rst,matrix_A[7742],matrix_B[142],mul_res1[7742]);
multi_7x28 multi_7x28_mod_7743(clk,rst,matrix_A[7743],matrix_B[143],mul_res1[7743]);
multi_7x28 multi_7x28_mod_7744(clk,rst,matrix_A[7744],matrix_B[144],mul_res1[7744]);
multi_7x28 multi_7x28_mod_7745(clk,rst,matrix_A[7745],matrix_B[145],mul_res1[7745]);
multi_7x28 multi_7x28_mod_7746(clk,rst,matrix_A[7746],matrix_B[146],mul_res1[7746]);
multi_7x28 multi_7x28_mod_7747(clk,rst,matrix_A[7747],matrix_B[147],mul_res1[7747]);
multi_7x28 multi_7x28_mod_7748(clk,rst,matrix_A[7748],matrix_B[148],mul_res1[7748]);
multi_7x28 multi_7x28_mod_7749(clk,rst,matrix_A[7749],matrix_B[149],mul_res1[7749]);
multi_7x28 multi_7x28_mod_7750(clk,rst,matrix_A[7750],matrix_B[150],mul_res1[7750]);
multi_7x28 multi_7x28_mod_7751(clk,rst,matrix_A[7751],matrix_B[151],mul_res1[7751]);
multi_7x28 multi_7x28_mod_7752(clk,rst,matrix_A[7752],matrix_B[152],mul_res1[7752]);
multi_7x28 multi_7x28_mod_7753(clk,rst,matrix_A[7753],matrix_B[153],mul_res1[7753]);
multi_7x28 multi_7x28_mod_7754(clk,rst,matrix_A[7754],matrix_B[154],mul_res1[7754]);
multi_7x28 multi_7x28_mod_7755(clk,rst,matrix_A[7755],matrix_B[155],mul_res1[7755]);
multi_7x28 multi_7x28_mod_7756(clk,rst,matrix_A[7756],matrix_B[156],mul_res1[7756]);
multi_7x28 multi_7x28_mod_7757(clk,rst,matrix_A[7757],matrix_B[157],mul_res1[7757]);
multi_7x28 multi_7x28_mod_7758(clk,rst,matrix_A[7758],matrix_B[158],mul_res1[7758]);
multi_7x28 multi_7x28_mod_7759(clk,rst,matrix_A[7759],matrix_B[159],mul_res1[7759]);
multi_7x28 multi_7x28_mod_7760(clk,rst,matrix_A[7760],matrix_B[160],mul_res1[7760]);
multi_7x28 multi_7x28_mod_7761(clk,rst,matrix_A[7761],matrix_B[161],mul_res1[7761]);
multi_7x28 multi_7x28_mod_7762(clk,rst,matrix_A[7762],matrix_B[162],mul_res1[7762]);
multi_7x28 multi_7x28_mod_7763(clk,rst,matrix_A[7763],matrix_B[163],mul_res1[7763]);
multi_7x28 multi_7x28_mod_7764(clk,rst,matrix_A[7764],matrix_B[164],mul_res1[7764]);
multi_7x28 multi_7x28_mod_7765(clk,rst,matrix_A[7765],matrix_B[165],mul_res1[7765]);
multi_7x28 multi_7x28_mod_7766(clk,rst,matrix_A[7766],matrix_B[166],mul_res1[7766]);
multi_7x28 multi_7x28_mod_7767(clk,rst,matrix_A[7767],matrix_B[167],mul_res1[7767]);
multi_7x28 multi_7x28_mod_7768(clk,rst,matrix_A[7768],matrix_B[168],mul_res1[7768]);
multi_7x28 multi_7x28_mod_7769(clk,rst,matrix_A[7769],matrix_B[169],mul_res1[7769]);
multi_7x28 multi_7x28_mod_7770(clk,rst,matrix_A[7770],matrix_B[170],mul_res1[7770]);
multi_7x28 multi_7x28_mod_7771(clk,rst,matrix_A[7771],matrix_B[171],mul_res1[7771]);
multi_7x28 multi_7x28_mod_7772(clk,rst,matrix_A[7772],matrix_B[172],mul_res1[7772]);
multi_7x28 multi_7x28_mod_7773(clk,rst,matrix_A[7773],matrix_B[173],mul_res1[7773]);
multi_7x28 multi_7x28_mod_7774(clk,rst,matrix_A[7774],matrix_B[174],mul_res1[7774]);
multi_7x28 multi_7x28_mod_7775(clk,rst,matrix_A[7775],matrix_B[175],mul_res1[7775]);
multi_7x28 multi_7x28_mod_7776(clk,rst,matrix_A[7776],matrix_B[176],mul_res1[7776]);
multi_7x28 multi_7x28_mod_7777(clk,rst,matrix_A[7777],matrix_B[177],mul_res1[7777]);
multi_7x28 multi_7x28_mod_7778(clk,rst,matrix_A[7778],matrix_B[178],mul_res1[7778]);
multi_7x28 multi_7x28_mod_7779(clk,rst,matrix_A[7779],matrix_B[179],mul_res1[7779]);
multi_7x28 multi_7x28_mod_7780(clk,rst,matrix_A[7780],matrix_B[180],mul_res1[7780]);
multi_7x28 multi_7x28_mod_7781(clk,rst,matrix_A[7781],matrix_B[181],mul_res1[7781]);
multi_7x28 multi_7x28_mod_7782(clk,rst,matrix_A[7782],matrix_B[182],mul_res1[7782]);
multi_7x28 multi_7x28_mod_7783(clk,rst,matrix_A[7783],matrix_B[183],mul_res1[7783]);
multi_7x28 multi_7x28_mod_7784(clk,rst,matrix_A[7784],matrix_B[184],mul_res1[7784]);
multi_7x28 multi_7x28_mod_7785(clk,rst,matrix_A[7785],matrix_B[185],mul_res1[7785]);
multi_7x28 multi_7x28_mod_7786(clk,rst,matrix_A[7786],matrix_B[186],mul_res1[7786]);
multi_7x28 multi_7x28_mod_7787(clk,rst,matrix_A[7787],matrix_B[187],mul_res1[7787]);
multi_7x28 multi_7x28_mod_7788(clk,rst,matrix_A[7788],matrix_B[188],mul_res1[7788]);
multi_7x28 multi_7x28_mod_7789(clk,rst,matrix_A[7789],matrix_B[189],mul_res1[7789]);
multi_7x28 multi_7x28_mod_7790(clk,rst,matrix_A[7790],matrix_B[190],mul_res1[7790]);
multi_7x28 multi_7x28_mod_7791(clk,rst,matrix_A[7791],matrix_B[191],mul_res1[7791]);
multi_7x28 multi_7x28_mod_7792(clk,rst,matrix_A[7792],matrix_B[192],mul_res1[7792]);
multi_7x28 multi_7x28_mod_7793(clk,rst,matrix_A[7793],matrix_B[193],mul_res1[7793]);
multi_7x28 multi_7x28_mod_7794(clk,rst,matrix_A[7794],matrix_B[194],mul_res1[7794]);
multi_7x28 multi_7x28_mod_7795(clk,rst,matrix_A[7795],matrix_B[195],mul_res1[7795]);
multi_7x28 multi_7x28_mod_7796(clk,rst,matrix_A[7796],matrix_B[196],mul_res1[7796]);
multi_7x28 multi_7x28_mod_7797(clk,rst,matrix_A[7797],matrix_B[197],mul_res1[7797]);
multi_7x28 multi_7x28_mod_7798(clk,rst,matrix_A[7798],matrix_B[198],mul_res1[7798]);
multi_7x28 multi_7x28_mod_7799(clk,rst,matrix_A[7799],matrix_B[199],mul_res1[7799]);
multi_7x28 multi_7x28_mod_7800(clk,rst,matrix_A[7800],matrix_B[0],mul_res1[7800]);
multi_7x28 multi_7x28_mod_7801(clk,rst,matrix_A[7801],matrix_B[1],mul_res1[7801]);
multi_7x28 multi_7x28_mod_7802(clk,rst,matrix_A[7802],matrix_B[2],mul_res1[7802]);
multi_7x28 multi_7x28_mod_7803(clk,rst,matrix_A[7803],matrix_B[3],mul_res1[7803]);
multi_7x28 multi_7x28_mod_7804(clk,rst,matrix_A[7804],matrix_B[4],mul_res1[7804]);
multi_7x28 multi_7x28_mod_7805(clk,rst,matrix_A[7805],matrix_B[5],mul_res1[7805]);
multi_7x28 multi_7x28_mod_7806(clk,rst,matrix_A[7806],matrix_B[6],mul_res1[7806]);
multi_7x28 multi_7x28_mod_7807(clk,rst,matrix_A[7807],matrix_B[7],mul_res1[7807]);
multi_7x28 multi_7x28_mod_7808(clk,rst,matrix_A[7808],matrix_B[8],mul_res1[7808]);
multi_7x28 multi_7x28_mod_7809(clk,rst,matrix_A[7809],matrix_B[9],mul_res1[7809]);
multi_7x28 multi_7x28_mod_7810(clk,rst,matrix_A[7810],matrix_B[10],mul_res1[7810]);
multi_7x28 multi_7x28_mod_7811(clk,rst,matrix_A[7811],matrix_B[11],mul_res1[7811]);
multi_7x28 multi_7x28_mod_7812(clk,rst,matrix_A[7812],matrix_B[12],mul_res1[7812]);
multi_7x28 multi_7x28_mod_7813(clk,rst,matrix_A[7813],matrix_B[13],mul_res1[7813]);
multi_7x28 multi_7x28_mod_7814(clk,rst,matrix_A[7814],matrix_B[14],mul_res1[7814]);
multi_7x28 multi_7x28_mod_7815(clk,rst,matrix_A[7815],matrix_B[15],mul_res1[7815]);
multi_7x28 multi_7x28_mod_7816(clk,rst,matrix_A[7816],matrix_B[16],mul_res1[7816]);
multi_7x28 multi_7x28_mod_7817(clk,rst,matrix_A[7817],matrix_B[17],mul_res1[7817]);
multi_7x28 multi_7x28_mod_7818(clk,rst,matrix_A[7818],matrix_B[18],mul_res1[7818]);
multi_7x28 multi_7x28_mod_7819(clk,rst,matrix_A[7819],matrix_B[19],mul_res1[7819]);
multi_7x28 multi_7x28_mod_7820(clk,rst,matrix_A[7820],matrix_B[20],mul_res1[7820]);
multi_7x28 multi_7x28_mod_7821(clk,rst,matrix_A[7821],matrix_B[21],mul_res1[7821]);
multi_7x28 multi_7x28_mod_7822(clk,rst,matrix_A[7822],matrix_B[22],mul_res1[7822]);
multi_7x28 multi_7x28_mod_7823(clk,rst,matrix_A[7823],matrix_B[23],mul_res1[7823]);
multi_7x28 multi_7x28_mod_7824(clk,rst,matrix_A[7824],matrix_B[24],mul_res1[7824]);
multi_7x28 multi_7x28_mod_7825(clk,rst,matrix_A[7825],matrix_B[25],mul_res1[7825]);
multi_7x28 multi_7x28_mod_7826(clk,rst,matrix_A[7826],matrix_B[26],mul_res1[7826]);
multi_7x28 multi_7x28_mod_7827(clk,rst,matrix_A[7827],matrix_B[27],mul_res1[7827]);
multi_7x28 multi_7x28_mod_7828(clk,rst,matrix_A[7828],matrix_B[28],mul_res1[7828]);
multi_7x28 multi_7x28_mod_7829(clk,rst,matrix_A[7829],matrix_B[29],mul_res1[7829]);
multi_7x28 multi_7x28_mod_7830(clk,rst,matrix_A[7830],matrix_B[30],mul_res1[7830]);
multi_7x28 multi_7x28_mod_7831(clk,rst,matrix_A[7831],matrix_B[31],mul_res1[7831]);
multi_7x28 multi_7x28_mod_7832(clk,rst,matrix_A[7832],matrix_B[32],mul_res1[7832]);
multi_7x28 multi_7x28_mod_7833(clk,rst,matrix_A[7833],matrix_B[33],mul_res1[7833]);
multi_7x28 multi_7x28_mod_7834(clk,rst,matrix_A[7834],matrix_B[34],mul_res1[7834]);
multi_7x28 multi_7x28_mod_7835(clk,rst,matrix_A[7835],matrix_B[35],mul_res1[7835]);
multi_7x28 multi_7x28_mod_7836(clk,rst,matrix_A[7836],matrix_B[36],mul_res1[7836]);
multi_7x28 multi_7x28_mod_7837(clk,rst,matrix_A[7837],matrix_B[37],mul_res1[7837]);
multi_7x28 multi_7x28_mod_7838(clk,rst,matrix_A[7838],matrix_B[38],mul_res1[7838]);
multi_7x28 multi_7x28_mod_7839(clk,rst,matrix_A[7839],matrix_B[39],mul_res1[7839]);
multi_7x28 multi_7x28_mod_7840(clk,rst,matrix_A[7840],matrix_B[40],mul_res1[7840]);
multi_7x28 multi_7x28_mod_7841(clk,rst,matrix_A[7841],matrix_B[41],mul_res1[7841]);
multi_7x28 multi_7x28_mod_7842(clk,rst,matrix_A[7842],matrix_B[42],mul_res1[7842]);
multi_7x28 multi_7x28_mod_7843(clk,rst,matrix_A[7843],matrix_B[43],mul_res1[7843]);
multi_7x28 multi_7x28_mod_7844(clk,rst,matrix_A[7844],matrix_B[44],mul_res1[7844]);
multi_7x28 multi_7x28_mod_7845(clk,rst,matrix_A[7845],matrix_B[45],mul_res1[7845]);
multi_7x28 multi_7x28_mod_7846(clk,rst,matrix_A[7846],matrix_B[46],mul_res1[7846]);
multi_7x28 multi_7x28_mod_7847(clk,rst,matrix_A[7847],matrix_B[47],mul_res1[7847]);
multi_7x28 multi_7x28_mod_7848(clk,rst,matrix_A[7848],matrix_B[48],mul_res1[7848]);
multi_7x28 multi_7x28_mod_7849(clk,rst,matrix_A[7849],matrix_B[49],mul_res1[7849]);
multi_7x28 multi_7x28_mod_7850(clk,rst,matrix_A[7850],matrix_B[50],mul_res1[7850]);
multi_7x28 multi_7x28_mod_7851(clk,rst,matrix_A[7851],matrix_B[51],mul_res1[7851]);
multi_7x28 multi_7x28_mod_7852(clk,rst,matrix_A[7852],matrix_B[52],mul_res1[7852]);
multi_7x28 multi_7x28_mod_7853(clk,rst,matrix_A[7853],matrix_B[53],mul_res1[7853]);
multi_7x28 multi_7x28_mod_7854(clk,rst,matrix_A[7854],matrix_B[54],mul_res1[7854]);
multi_7x28 multi_7x28_mod_7855(clk,rst,matrix_A[7855],matrix_B[55],mul_res1[7855]);
multi_7x28 multi_7x28_mod_7856(clk,rst,matrix_A[7856],matrix_B[56],mul_res1[7856]);
multi_7x28 multi_7x28_mod_7857(clk,rst,matrix_A[7857],matrix_B[57],mul_res1[7857]);
multi_7x28 multi_7x28_mod_7858(clk,rst,matrix_A[7858],matrix_B[58],mul_res1[7858]);
multi_7x28 multi_7x28_mod_7859(clk,rst,matrix_A[7859],matrix_B[59],mul_res1[7859]);
multi_7x28 multi_7x28_mod_7860(clk,rst,matrix_A[7860],matrix_B[60],mul_res1[7860]);
multi_7x28 multi_7x28_mod_7861(clk,rst,matrix_A[7861],matrix_B[61],mul_res1[7861]);
multi_7x28 multi_7x28_mod_7862(clk,rst,matrix_A[7862],matrix_B[62],mul_res1[7862]);
multi_7x28 multi_7x28_mod_7863(clk,rst,matrix_A[7863],matrix_B[63],mul_res1[7863]);
multi_7x28 multi_7x28_mod_7864(clk,rst,matrix_A[7864],matrix_B[64],mul_res1[7864]);
multi_7x28 multi_7x28_mod_7865(clk,rst,matrix_A[7865],matrix_B[65],mul_res1[7865]);
multi_7x28 multi_7x28_mod_7866(clk,rst,matrix_A[7866],matrix_B[66],mul_res1[7866]);
multi_7x28 multi_7x28_mod_7867(clk,rst,matrix_A[7867],matrix_B[67],mul_res1[7867]);
multi_7x28 multi_7x28_mod_7868(clk,rst,matrix_A[7868],matrix_B[68],mul_res1[7868]);
multi_7x28 multi_7x28_mod_7869(clk,rst,matrix_A[7869],matrix_B[69],mul_res1[7869]);
multi_7x28 multi_7x28_mod_7870(clk,rst,matrix_A[7870],matrix_B[70],mul_res1[7870]);
multi_7x28 multi_7x28_mod_7871(clk,rst,matrix_A[7871],matrix_B[71],mul_res1[7871]);
multi_7x28 multi_7x28_mod_7872(clk,rst,matrix_A[7872],matrix_B[72],mul_res1[7872]);
multi_7x28 multi_7x28_mod_7873(clk,rst,matrix_A[7873],matrix_B[73],mul_res1[7873]);
multi_7x28 multi_7x28_mod_7874(clk,rst,matrix_A[7874],matrix_B[74],mul_res1[7874]);
multi_7x28 multi_7x28_mod_7875(clk,rst,matrix_A[7875],matrix_B[75],mul_res1[7875]);
multi_7x28 multi_7x28_mod_7876(clk,rst,matrix_A[7876],matrix_B[76],mul_res1[7876]);
multi_7x28 multi_7x28_mod_7877(clk,rst,matrix_A[7877],matrix_B[77],mul_res1[7877]);
multi_7x28 multi_7x28_mod_7878(clk,rst,matrix_A[7878],matrix_B[78],mul_res1[7878]);
multi_7x28 multi_7x28_mod_7879(clk,rst,matrix_A[7879],matrix_B[79],mul_res1[7879]);
multi_7x28 multi_7x28_mod_7880(clk,rst,matrix_A[7880],matrix_B[80],mul_res1[7880]);
multi_7x28 multi_7x28_mod_7881(clk,rst,matrix_A[7881],matrix_B[81],mul_res1[7881]);
multi_7x28 multi_7x28_mod_7882(clk,rst,matrix_A[7882],matrix_B[82],mul_res1[7882]);
multi_7x28 multi_7x28_mod_7883(clk,rst,matrix_A[7883],matrix_B[83],mul_res1[7883]);
multi_7x28 multi_7x28_mod_7884(clk,rst,matrix_A[7884],matrix_B[84],mul_res1[7884]);
multi_7x28 multi_7x28_mod_7885(clk,rst,matrix_A[7885],matrix_B[85],mul_res1[7885]);
multi_7x28 multi_7x28_mod_7886(clk,rst,matrix_A[7886],matrix_B[86],mul_res1[7886]);
multi_7x28 multi_7x28_mod_7887(clk,rst,matrix_A[7887],matrix_B[87],mul_res1[7887]);
multi_7x28 multi_7x28_mod_7888(clk,rst,matrix_A[7888],matrix_B[88],mul_res1[7888]);
multi_7x28 multi_7x28_mod_7889(clk,rst,matrix_A[7889],matrix_B[89],mul_res1[7889]);
multi_7x28 multi_7x28_mod_7890(clk,rst,matrix_A[7890],matrix_B[90],mul_res1[7890]);
multi_7x28 multi_7x28_mod_7891(clk,rst,matrix_A[7891],matrix_B[91],mul_res1[7891]);
multi_7x28 multi_7x28_mod_7892(clk,rst,matrix_A[7892],matrix_B[92],mul_res1[7892]);
multi_7x28 multi_7x28_mod_7893(clk,rst,matrix_A[7893],matrix_B[93],mul_res1[7893]);
multi_7x28 multi_7x28_mod_7894(clk,rst,matrix_A[7894],matrix_B[94],mul_res1[7894]);
multi_7x28 multi_7x28_mod_7895(clk,rst,matrix_A[7895],matrix_B[95],mul_res1[7895]);
multi_7x28 multi_7x28_mod_7896(clk,rst,matrix_A[7896],matrix_B[96],mul_res1[7896]);
multi_7x28 multi_7x28_mod_7897(clk,rst,matrix_A[7897],matrix_B[97],mul_res1[7897]);
multi_7x28 multi_7x28_mod_7898(clk,rst,matrix_A[7898],matrix_B[98],mul_res1[7898]);
multi_7x28 multi_7x28_mod_7899(clk,rst,matrix_A[7899],matrix_B[99],mul_res1[7899]);
multi_7x28 multi_7x28_mod_7900(clk,rst,matrix_A[7900],matrix_B[100],mul_res1[7900]);
multi_7x28 multi_7x28_mod_7901(clk,rst,matrix_A[7901],matrix_B[101],mul_res1[7901]);
multi_7x28 multi_7x28_mod_7902(clk,rst,matrix_A[7902],matrix_B[102],mul_res1[7902]);
multi_7x28 multi_7x28_mod_7903(clk,rst,matrix_A[7903],matrix_B[103],mul_res1[7903]);
multi_7x28 multi_7x28_mod_7904(clk,rst,matrix_A[7904],matrix_B[104],mul_res1[7904]);
multi_7x28 multi_7x28_mod_7905(clk,rst,matrix_A[7905],matrix_B[105],mul_res1[7905]);
multi_7x28 multi_7x28_mod_7906(clk,rst,matrix_A[7906],matrix_B[106],mul_res1[7906]);
multi_7x28 multi_7x28_mod_7907(clk,rst,matrix_A[7907],matrix_B[107],mul_res1[7907]);
multi_7x28 multi_7x28_mod_7908(clk,rst,matrix_A[7908],matrix_B[108],mul_res1[7908]);
multi_7x28 multi_7x28_mod_7909(clk,rst,matrix_A[7909],matrix_B[109],mul_res1[7909]);
multi_7x28 multi_7x28_mod_7910(clk,rst,matrix_A[7910],matrix_B[110],mul_res1[7910]);
multi_7x28 multi_7x28_mod_7911(clk,rst,matrix_A[7911],matrix_B[111],mul_res1[7911]);
multi_7x28 multi_7x28_mod_7912(clk,rst,matrix_A[7912],matrix_B[112],mul_res1[7912]);
multi_7x28 multi_7x28_mod_7913(clk,rst,matrix_A[7913],matrix_B[113],mul_res1[7913]);
multi_7x28 multi_7x28_mod_7914(clk,rst,matrix_A[7914],matrix_B[114],mul_res1[7914]);
multi_7x28 multi_7x28_mod_7915(clk,rst,matrix_A[7915],matrix_B[115],mul_res1[7915]);
multi_7x28 multi_7x28_mod_7916(clk,rst,matrix_A[7916],matrix_B[116],mul_res1[7916]);
multi_7x28 multi_7x28_mod_7917(clk,rst,matrix_A[7917],matrix_B[117],mul_res1[7917]);
multi_7x28 multi_7x28_mod_7918(clk,rst,matrix_A[7918],matrix_B[118],mul_res1[7918]);
multi_7x28 multi_7x28_mod_7919(clk,rst,matrix_A[7919],matrix_B[119],mul_res1[7919]);
multi_7x28 multi_7x28_mod_7920(clk,rst,matrix_A[7920],matrix_B[120],mul_res1[7920]);
multi_7x28 multi_7x28_mod_7921(clk,rst,matrix_A[7921],matrix_B[121],mul_res1[7921]);
multi_7x28 multi_7x28_mod_7922(clk,rst,matrix_A[7922],matrix_B[122],mul_res1[7922]);
multi_7x28 multi_7x28_mod_7923(clk,rst,matrix_A[7923],matrix_B[123],mul_res1[7923]);
multi_7x28 multi_7x28_mod_7924(clk,rst,matrix_A[7924],matrix_B[124],mul_res1[7924]);
multi_7x28 multi_7x28_mod_7925(clk,rst,matrix_A[7925],matrix_B[125],mul_res1[7925]);
multi_7x28 multi_7x28_mod_7926(clk,rst,matrix_A[7926],matrix_B[126],mul_res1[7926]);
multi_7x28 multi_7x28_mod_7927(clk,rst,matrix_A[7927],matrix_B[127],mul_res1[7927]);
multi_7x28 multi_7x28_mod_7928(clk,rst,matrix_A[7928],matrix_B[128],mul_res1[7928]);
multi_7x28 multi_7x28_mod_7929(clk,rst,matrix_A[7929],matrix_B[129],mul_res1[7929]);
multi_7x28 multi_7x28_mod_7930(clk,rst,matrix_A[7930],matrix_B[130],mul_res1[7930]);
multi_7x28 multi_7x28_mod_7931(clk,rst,matrix_A[7931],matrix_B[131],mul_res1[7931]);
multi_7x28 multi_7x28_mod_7932(clk,rst,matrix_A[7932],matrix_B[132],mul_res1[7932]);
multi_7x28 multi_7x28_mod_7933(clk,rst,matrix_A[7933],matrix_B[133],mul_res1[7933]);
multi_7x28 multi_7x28_mod_7934(clk,rst,matrix_A[7934],matrix_B[134],mul_res1[7934]);
multi_7x28 multi_7x28_mod_7935(clk,rst,matrix_A[7935],matrix_B[135],mul_res1[7935]);
multi_7x28 multi_7x28_mod_7936(clk,rst,matrix_A[7936],matrix_B[136],mul_res1[7936]);
multi_7x28 multi_7x28_mod_7937(clk,rst,matrix_A[7937],matrix_B[137],mul_res1[7937]);
multi_7x28 multi_7x28_mod_7938(clk,rst,matrix_A[7938],matrix_B[138],mul_res1[7938]);
multi_7x28 multi_7x28_mod_7939(clk,rst,matrix_A[7939],matrix_B[139],mul_res1[7939]);
multi_7x28 multi_7x28_mod_7940(clk,rst,matrix_A[7940],matrix_B[140],mul_res1[7940]);
multi_7x28 multi_7x28_mod_7941(clk,rst,matrix_A[7941],matrix_B[141],mul_res1[7941]);
multi_7x28 multi_7x28_mod_7942(clk,rst,matrix_A[7942],matrix_B[142],mul_res1[7942]);
multi_7x28 multi_7x28_mod_7943(clk,rst,matrix_A[7943],matrix_B[143],mul_res1[7943]);
multi_7x28 multi_7x28_mod_7944(clk,rst,matrix_A[7944],matrix_B[144],mul_res1[7944]);
multi_7x28 multi_7x28_mod_7945(clk,rst,matrix_A[7945],matrix_B[145],mul_res1[7945]);
multi_7x28 multi_7x28_mod_7946(clk,rst,matrix_A[7946],matrix_B[146],mul_res1[7946]);
multi_7x28 multi_7x28_mod_7947(clk,rst,matrix_A[7947],matrix_B[147],mul_res1[7947]);
multi_7x28 multi_7x28_mod_7948(clk,rst,matrix_A[7948],matrix_B[148],mul_res1[7948]);
multi_7x28 multi_7x28_mod_7949(clk,rst,matrix_A[7949],matrix_B[149],mul_res1[7949]);
multi_7x28 multi_7x28_mod_7950(clk,rst,matrix_A[7950],matrix_B[150],mul_res1[7950]);
multi_7x28 multi_7x28_mod_7951(clk,rst,matrix_A[7951],matrix_B[151],mul_res1[7951]);
multi_7x28 multi_7x28_mod_7952(clk,rst,matrix_A[7952],matrix_B[152],mul_res1[7952]);
multi_7x28 multi_7x28_mod_7953(clk,rst,matrix_A[7953],matrix_B[153],mul_res1[7953]);
multi_7x28 multi_7x28_mod_7954(clk,rst,matrix_A[7954],matrix_B[154],mul_res1[7954]);
multi_7x28 multi_7x28_mod_7955(clk,rst,matrix_A[7955],matrix_B[155],mul_res1[7955]);
multi_7x28 multi_7x28_mod_7956(clk,rst,matrix_A[7956],matrix_B[156],mul_res1[7956]);
multi_7x28 multi_7x28_mod_7957(clk,rst,matrix_A[7957],matrix_B[157],mul_res1[7957]);
multi_7x28 multi_7x28_mod_7958(clk,rst,matrix_A[7958],matrix_B[158],mul_res1[7958]);
multi_7x28 multi_7x28_mod_7959(clk,rst,matrix_A[7959],matrix_B[159],mul_res1[7959]);
multi_7x28 multi_7x28_mod_7960(clk,rst,matrix_A[7960],matrix_B[160],mul_res1[7960]);
multi_7x28 multi_7x28_mod_7961(clk,rst,matrix_A[7961],matrix_B[161],mul_res1[7961]);
multi_7x28 multi_7x28_mod_7962(clk,rst,matrix_A[7962],matrix_B[162],mul_res1[7962]);
multi_7x28 multi_7x28_mod_7963(clk,rst,matrix_A[7963],matrix_B[163],mul_res1[7963]);
multi_7x28 multi_7x28_mod_7964(clk,rst,matrix_A[7964],matrix_B[164],mul_res1[7964]);
multi_7x28 multi_7x28_mod_7965(clk,rst,matrix_A[7965],matrix_B[165],mul_res1[7965]);
multi_7x28 multi_7x28_mod_7966(clk,rst,matrix_A[7966],matrix_B[166],mul_res1[7966]);
multi_7x28 multi_7x28_mod_7967(clk,rst,matrix_A[7967],matrix_B[167],mul_res1[7967]);
multi_7x28 multi_7x28_mod_7968(clk,rst,matrix_A[7968],matrix_B[168],mul_res1[7968]);
multi_7x28 multi_7x28_mod_7969(clk,rst,matrix_A[7969],matrix_B[169],mul_res1[7969]);
multi_7x28 multi_7x28_mod_7970(clk,rst,matrix_A[7970],matrix_B[170],mul_res1[7970]);
multi_7x28 multi_7x28_mod_7971(clk,rst,matrix_A[7971],matrix_B[171],mul_res1[7971]);
multi_7x28 multi_7x28_mod_7972(clk,rst,matrix_A[7972],matrix_B[172],mul_res1[7972]);
multi_7x28 multi_7x28_mod_7973(clk,rst,matrix_A[7973],matrix_B[173],mul_res1[7973]);
multi_7x28 multi_7x28_mod_7974(clk,rst,matrix_A[7974],matrix_B[174],mul_res1[7974]);
multi_7x28 multi_7x28_mod_7975(clk,rst,matrix_A[7975],matrix_B[175],mul_res1[7975]);
multi_7x28 multi_7x28_mod_7976(clk,rst,matrix_A[7976],matrix_B[176],mul_res1[7976]);
multi_7x28 multi_7x28_mod_7977(clk,rst,matrix_A[7977],matrix_B[177],mul_res1[7977]);
multi_7x28 multi_7x28_mod_7978(clk,rst,matrix_A[7978],matrix_B[178],mul_res1[7978]);
multi_7x28 multi_7x28_mod_7979(clk,rst,matrix_A[7979],matrix_B[179],mul_res1[7979]);
multi_7x28 multi_7x28_mod_7980(clk,rst,matrix_A[7980],matrix_B[180],mul_res1[7980]);
multi_7x28 multi_7x28_mod_7981(clk,rst,matrix_A[7981],matrix_B[181],mul_res1[7981]);
multi_7x28 multi_7x28_mod_7982(clk,rst,matrix_A[7982],matrix_B[182],mul_res1[7982]);
multi_7x28 multi_7x28_mod_7983(clk,rst,matrix_A[7983],matrix_B[183],mul_res1[7983]);
multi_7x28 multi_7x28_mod_7984(clk,rst,matrix_A[7984],matrix_B[184],mul_res1[7984]);
multi_7x28 multi_7x28_mod_7985(clk,rst,matrix_A[7985],matrix_B[185],mul_res1[7985]);
multi_7x28 multi_7x28_mod_7986(clk,rst,matrix_A[7986],matrix_B[186],mul_res1[7986]);
multi_7x28 multi_7x28_mod_7987(clk,rst,matrix_A[7987],matrix_B[187],mul_res1[7987]);
multi_7x28 multi_7x28_mod_7988(clk,rst,matrix_A[7988],matrix_B[188],mul_res1[7988]);
multi_7x28 multi_7x28_mod_7989(clk,rst,matrix_A[7989],matrix_B[189],mul_res1[7989]);
multi_7x28 multi_7x28_mod_7990(clk,rst,matrix_A[7990],matrix_B[190],mul_res1[7990]);
multi_7x28 multi_7x28_mod_7991(clk,rst,matrix_A[7991],matrix_B[191],mul_res1[7991]);
multi_7x28 multi_7x28_mod_7992(clk,rst,matrix_A[7992],matrix_B[192],mul_res1[7992]);
multi_7x28 multi_7x28_mod_7993(clk,rst,matrix_A[7993],matrix_B[193],mul_res1[7993]);
multi_7x28 multi_7x28_mod_7994(clk,rst,matrix_A[7994],matrix_B[194],mul_res1[7994]);
multi_7x28 multi_7x28_mod_7995(clk,rst,matrix_A[7995],matrix_B[195],mul_res1[7995]);
multi_7x28 multi_7x28_mod_7996(clk,rst,matrix_A[7996],matrix_B[196],mul_res1[7996]);
multi_7x28 multi_7x28_mod_7997(clk,rst,matrix_A[7997],matrix_B[197],mul_res1[7997]);
multi_7x28 multi_7x28_mod_7998(clk,rst,matrix_A[7998],matrix_B[198],mul_res1[7998]);
multi_7x28 multi_7x28_mod_7999(clk,rst,matrix_A[7999],matrix_B[199],mul_res1[7999]);
multi_7x28 multi_7x28_mod_8000(clk,rst,matrix_A[8000],matrix_B[0],mul_res1[8000]);
multi_7x28 multi_7x28_mod_8001(clk,rst,matrix_A[8001],matrix_B[1],mul_res1[8001]);
multi_7x28 multi_7x28_mod_8002(clk,rst,matrix_A[8002],matrix_B[2],mul_res1[8002]);
multi_7x28 multi_7x28_mod_8003(clk,rst,matrix_A[8003],matrix_B[3],mul_res1[8003]);
multi_7x28 multi_7x28_mod_8004(clk,rst,matrix_A[8004],matrix_B[4],mul_res1[8004]);
multi_7x28 multi_7x28_mod_8005(clk,rst,matrix_A[8005],matrix_B[5],mul_res1[8005]);
multi_7x28 multi_7x28_mod_8006(clk,rst,matrix_A[8006],matrix_B[6],mul_res1[8006]);
multi_7x28 multi_7x28_mod_8007(clk,rst,matrix_A[8007],matrix_B[7],mul_res1[8007]);
multi_7x28 multi_7x28_mod_8008(clk,rst,matrix_A[8008],matrix_B[8],mul_res1[8008]);
multi_7x28 multi_7x28_mod_8009(clk,rst,matrix_A[8009],matrix_B[9],mul_res1[8009]);
multi_7x28 multi_7x28_mod_8010(clk,rst,matrix_A[8010],matrix_B[10],mul_res1[8010]);
multi_7x28 multi_7x28_mod_8011(clk,rst,matrix_A[8011],matrix_B[11],mul_res1[8011]);
multi_7x28 multi_7x28_mod_8012(clk,rst,matrix_A[8012],matrix_B[12],mul_res1[8012]);
multi_7x28 multi_7x28_mod_8013(clk,rst,matrix_A[8013],matrix_B[13],mul_res1[8013]);
multi_7x28 multi_7x28_mod_8014(clk,rst,matrix_A[8014],matrix_B[14],mul_res1[8014]);
multi_7x28 multi_7x28_mod_8015(clk,rst,matrix_A[8015],matrix_B[15],mul_res1[8015]);
multi_7x28 multi_7x28_mod_8016(clk,rst,matrix_A[8016],matrix_B[16],mul_res1[8016]);
multi_7x28 multi_7x28_mod_8017(clk,rst,matrix_A[8017],matrix_B[17],mul_res1[8017]);
multi_7x28 multi_7x28_mod_8018(clk,rst,matrix_A[8018],matrix_B[18],mul_res1[8018]);
multi_7x28 multi_7x28_mod_8019(clk,rst,matrix_A[8019],matrix_B[19],mul_res1[8019]);
multi_7x28 multi_7x28_mod_8020(clk,rst,matrix_A[8020],matrix_B[20],mul_res1[8020]);
multi_7x28 multi_7x28_mod_8021(clk,rst,matrix_A[8021],matrix_B[21],mul_res1[8021]);
multi_7x28 multi_7x28_mod_8022(clk,rst,matrix_A[8022],matrix_B[22],mul_res1[8022]);
multi_7x28 multi_7x28_mod_8023(clk,rst,matrix_A[8023],matrix_B[23],mul_res1[8023]);
multi_7x28 multi_7x28_mod_8024(clk,rst,matrix_A[8024],matrix_B[24],mul_res1[8024]);
multi_7x28 multi_7x28_mod_8025(clk,rst,matrix_A[8025],matrix_B[25],mul_res1[8025]);
multi_7x28 multi_7x28_mod_8026(clk,rst,matrix_A[8026],matrix_B[26],mul_res1[8026]);
multi_7x28 multi_7x28_mod_8027(clk,rst,matrix_A[8027],matrix_B[27],mul_res1[8027]);
multi_7x28 multi_7x28_mod_8028(clk,rst,matrix_A[8028],matrix_B[28],mul_res1[8028]);
multi_7x28 multi_7x28_mod_8029(clk,rst,matrix_A[8029],matrix_B[29],mul_res1[8029]);
multi_7x28 multi_7x28_mod_8030(clk,rst,matrix_A[8030],matrix_B[30],mul_res1[8030]);
multi_7x28 multi_7x28_mod_8031(clk,rst,matrix_A[8031],matrix_B[31],mul_res1[8031]);
multi_7x28 multi_7x28_mod_8032(clk,rst,matrix_A[8032],matrix_B[32],mul_res1[8032]);
multi_7x28 multi_7x28_mod_8033(clk,rst,matrix_A[8033],matrix_B[33],mul_res1[8033]);
multi_7x28 multi_7x28_mod_8034(clk,rst,matrix_A[8034],matrix_B[34],mul_res1[8034]);
multi_7x28 multi_7x28_mod_8035(clk,rst,matrix_A[8035],matrix_B[35],mul_res1[8035]);
multi_7x28 multi_7x28_mod_8036(clk,rst,matrix_A[8036],matrix_B[36],mul_res1[8036]);
multi_7x28 multi_7x28_mod_8037(clk,rst,matrix_A[8037],matrix_B[37],mul_res1[8037]);
multi_7x28 multi_7x28_mod_8038(clk,rst,matrix_A[8038],matrix_B[38],mul_res1[8038]);
multi_7x28 multi_7x28_mod_8039(clk,rst,matrix_A[8039],matrix_B[39],mul_res1[8039]);
multi_7x28 multi_7x28_mod_8040(clk,rst,matrix_A[8040],matrix_B[40],mul_res1[8040]);
multi_7x28 multi_7x28_mod_8041(clk,rst,matrix_A[8041],matrix_B[41],mul_res1[8041]);
multi_7x28 multi_7x28_mod_8042(clk,rst,matrix_A[8042],matrix_B[42],mul_res1[8042]);
multi_7x28 multi_7x28_mod_8043(clk,rst,matrix_A[8043],matrix_B[43],mul_res1[8043]);
multi_7x28 multi_7x28_mod_8044(clk,rst,matrix_A[8044],matrix_B[44],mul_res1[8044]);
multi_7x28 multi_7x28_mod_8045(clk,rst,matrix_A[8045],matrix_B[45],mul_res1[8045]);
multi_7x28 multi_7x28_mod_8046(clk,rst,matrix_A[8046],matrix_B[46],mul_res1[8046]);
multi_7x28 multi_7x28_mod_8047(clk,rst,matrix_A[8047],matrix_B[47],mul_res1[8047]);
multi_7x28 multi_7x28_mod_8048(clk,rst,matrix_A[8048],matrix_B[48],mul_res1[8048]);
multi_7x28 multi_7x28_mod_8049(clk,rst,matrix_A[8049],matrix_B[49],mul_res1[8049]);
multi_7x28 multi_7x28_mod_8050(clk,rst,matrix_A[8050],matrix_B[50],mul_res1[8050]);
multi_7x28 multi_7x28_mod_8051(clk,rst,matrix_A[8051],matrix_B[51],mul_res1[8051]);
multi_7x28 multi_7x28_mod_8052(clk,rst,matrix_A[8052],matrix_B[52],mul_res1[8052]);
multi_7x28 multi_7x28_mod_8053(clk,rst,matrix_A[8053],matrix_B[53],mul_res1[8053]);
multi_7x28 multi_7x28_mod_8054(clk,rst,matrix_A[8054],matrix_B[54],mul_res1[8054]);
multi_7x28 multi_7x28_mod_8055(clk,rst,matrix_A[8055],matrix_B[55],mul_res1[8055]);
multi_7x28 multi_7x28_mod_8056(clk,rst,matrix_A[8056],matrix_B[56],mul_res1[8056]);
multi_7x28 multi_7x28_mod_8057(clk,rst,matrix_A[8057],matrix_B[57],mul_res1[8057]);
multi_7x28 multi_7x28_mod_8058(clk,rst,matrix_A[8058],matrix_B[58],mul_res1[8058]);
multi_7x28 multi_7x28_mod_8059(clk,rst,matrix_A[8059],matrix_B[59],mul_res1[8059]);
multi_7x28 multi_7x28_mod_8060(clk,rst,matrix_A[8060],matrix_B[60],mul_res1[8060]);
multi_7x28 multi_7x28_mod_8061(clk,rst,matrix_A[8061],matrix_B[61],mul_res1[8061]);
multi_7x28 multi_7x28_mod_8062(clk,rst,matrix_A[8062],matrix_B[62],mul_res1[8062]);
multi_7x28 multi_7x28_mod_8063(clk,rst,matrix_A[8063],matrix_B[63],mul_res1[8063]);
multi_7x28 multi_7x28_mod_8064(clk,rst,matrix_A[8064],matrix_B[64],mul_res1[8064]);
multi_7x28 multi_7x28_mod_8065(clk,rst,matrix_A[8065],matrix_B[65],mul_res1[8065]);
multi_7x28 multi_7x28_mod_8066(clk,rst,matrix_A[8066],matrix_B[66],mul_res1[8066]);
multi_7x28 multi_7x28_mod_8067(clk,rst,matrix_A[8067],matrix_B[67],mul_res1[8067]);
multi_7x28 multi_7x28_mod_8068(clk,rst,matrix_A[8068],matrix_B[68],mul_res1[8068]);
multi_7x28 multi_7x28_mod_8069(clk,rst,matrix_A[8069],matrix_B[69],mul_res1[8069]);
multi_7x28 multi_7x28_mod_8070(clk,rst,matrix_A[8070],matrix_B[70],mul_res1[8070]);
multi_7x28 multi_7x28_mod_8071(clk,rst,matrix_A[8071],matrix_B[71],mul_res1[8071]);
multi_7x28 multi_7x28_mod_8072(clk,rst,matrix_A[8072],matrix_B[72],mul_res1[8072]);
multi_7x28 multi_7x28_mod_8073(clk,rst,matrix_A[8073],matrix_B[73],mul_res1[8073]);
multi_7x28 multi_7x28_mod_8074(clk,rst,matrix_A[8074],matrix_B[74],mul_res1[8074]);
multi_7x28 multi_7x28_mod_8075(clk,rst,matrix_A[8075],matrix_B[75],mul_res1[8075]);
multi_7x28 multi_7x28_mod_8076(clk,rst,matrix_A[8076],matrix_B[76],mul_res1[8076]);
multi_7x28 multi_7x28_mod_8077(clk,rst,matrix_A[8077],matrix_B[77],mul_res1[8077]);
multi_7x28 multi_7x28_mod_8078(clk,rst,matrix_A[8078],matrix_B[78],mul_res1[8078]);
multi_7x28 multi_7x28_mod_8079(clk,rst,matrix_A[8079],matrix_B[79],mul_res1[8079]);
multi_7x28 multi_7x28_mod_8080(clk,rst,matrix_A[8080],matrix_B[80],mul_res1[8080]);
multi_7x28 multi_7x28_mod_8081(clk,rst,matrix_A[8081],matrix_B[81],mul_res1[8081]);
multi_7x28 multi_7x28_mod_8082(clk,rst,matrix_A[8082],matrix_B[82],mul_res1[8082]);
multi_7x28 multi_7x28_mod_8083(clk,rst,matrix_A[8083],matrix_B[83],mul_res1[8083]);
multi_7x28 multi_7x28_mod_8084(clk,rst,matrix_A[8084],matrix_B[84],mul_res1[8084]);
multi_7x28 multi_7x28_mod_8085(clk,rst,matrix_A[8085],matrix_B[85],mul_res1[8085]);
multi_7x28 multi_7x28_mod_8086(clk,rst,matrix_A[8086],matrix_B[86],mul_res1[8086]);
multi_7x28 multi_7x28_mod_8087(clk,rst,matrix_A[8087],matrix_B[87],mul_res1[8087]);
multi_7x28 multi_7x28_mod_8088(clk,rst,matrix_A[8088],matrix_B[88],mul_res1[8088]);
multi_7x28 multi_7x28_mod_8089(clk,rst,matrix_A[8089],matrix_B[89],mul_res1[8089]);
multi_7x28 multi_7x28_mod_8090(clk,rst,matrix_A[8090],matrix_B[90],mul_res1[8090]);
multi_7x28 multi_7x28_mod_8091(clk,rst,matrix_A[8091],matrix_B[91],mul_res1[8091]);
multi_7x28 multi_7x28_mod_8092(clk,rst,matrix_A[8092],matrix_B[92],mul_res1[8092]);
multi_7x28 multi_7x28_mod_8093(clk,rst,matrix_A[8093],matrix_B[93],mul_res1[8093]);
multi_7x28 multi_7x28_mod_8094(clk,rst,matrix_A[8094],matrix_B[94],mul_res1[8094]);
multi_7x28 multi_7x28_mod_8095(clk,rst,matrix_A[8095],matrix_B[95],mul_res1[8095]);
multi_7x28 multi_7x28_mod_8096(clk,rst,matrix_A[8096],matrix_B[96],mul_res1[8096]);
multi_7x28 multi_7x28_mod_8097(clk,rst,matrix_A[8097],matrix_B[97],mul_res1[8097]);
multi_7x28 multi_7x28_mod_8098(clk,rst,matrix_A[8098],matrix_B[98],mul_res1[8098]);
multi_7x28 multi_7x28_mod_8099(clk,rst,matrix_A[8099],matrix_B[99],mul_res1[8099]);
multi_7x28 multi_7x28_mod_8100(clk,rst,matrix_A[8100],matrix_B[100],mul_res1[8100]);
multi_7x28 multi_7x28_mod_8101(clk,rst,matrix_A[8101],matrix_B[101],mul_res1[8101]);
multi_7x28 multi_7x28_mod_8102(clk,rst,matrix_A[8102],matrix_B[102],mul_res1[8102]);
multi_7x28 multi_7x28_mod_8103(clk,rst,matrix_A[8103],matrix_B[103],mul_res1[8103]);
multi_7x28 multi_7x28_mod_8104(clk,rst,matrix_A[8104],matrix_B[104],mul_res1[8104]);
multi_7x28 multi_7x28_mod_8105(clk,rst,matrix_A[8105],matrix_B[105],mul_res1[8105]);
multi_7x28 multi_7x28_mod_8106(clk,rst,matrix_A[8106],matrix_B[106],mul_res1[8106]);
multi_7x28 multi_7x28_mod_8107(clk,rst,matrix_A[8107],matrix_B[107],mul_res1[8107]);
multi_7x28 multi_7x28_mod_8108(clk,rst,matrix_A[8108],matrix_B[108],mul_res1[8108]);
multi_7x28 multi_7x28_mod_8109(clk,rst,matrix_A[8109],matrix_B[109],mul_res1[8109]);
multi_7x28 multi_7x28_mod_8110(clk,rst,matrix_A[8110],matrix_B[110],mul_res1[8110]);
multi_7x28 multi_7x28_mod_8111(clk,rst,matrix_A[8111],matrix_B[111],mul_res1[8111]);
multi_7x28 multi_7x28_mod_8112(clk,rst,matrix_A[8112],matrix_B[112],mul_res1[8112]);
multi_7x28 multi_7x28_mod_8113(clk,rst,matrix_A[8113],matrix_B[113],mul_res1[8113]);
multi_7x28 multi_7x28_mod_8114(clk,rst,matrix_A[8114],matrix_B[114],mul_res1[8114]);
multi_7x28 multi_7x28_mod_8115(clk,rst,matrix_A[8115],matrix_B[115],mul_res1[8115]);
multi_7x28 multi_7x28_mod_8116(clk,rst,matrix_A[8116],matrix_B[116],mul_res1[8116]);
multi_7x28 multi_7x28_mod_8117(clk,rst,matrix_A[8117],matrix_B[117],mul_res1[8117]);
multi_7x28 multi_7x28_mod_8118(clk,rst,matrix_A[8118],matrix_B[118],mul_res1[8118]);
multi_7x28 multi_7x28_mod_8119(clk,rst,matrix_A[8119],matrix_B[119],mul_res1[8119]);
multi_7x28 multi_7x28_mod_8120(clk,rst,matrix_A[8120],matrix_B[120],mul_res1[8120]);
multi_7x28 multi_7x28_mod_8121(clk,rst,matrix_A[8121],matrix_B[121],mul_res1[8121]);
multi_7x28 multi_7x28_mod_8122(clk,rst,matrix_A[8122],matrix_B[122],mul_res1[8122]);
multi_7x28 multi_7x28_mod_8123(clk,rst,matrix_A[8123],matrix_B[123],mul_res1[8123]);
multi_7x28 multi_7x28_mod_8124(clk,rst,matrix_A[8124],matrix_B[124],mul_res1[8124]);
multi_7x28 multi_7x28_mod_8125(clk,rst,matrix_A[8125],matrix_B[125],mul_res1[8125]);
multi_7x28 multi_7x28_mod_8126(clk,rst,matrix_A[8126],matrix_B[126],mul_res1[8126]);
multi_7x28 multi_7x28_mod_8127(clk,rst,matrix_A[8127],matrix_B[127],mul_res1[8127]);
multi_7x28 multi_7x28_mod_8128(clk,rst,matrix_A[8128],matrix_B[128],mul_res1[8128]);
multi_7x28 multi_7x28_mod_8129(clk,rst,matrix_A[8129],matrix_B[129],mul_res1[8129]);
multi_7x28 multi_7x28_mod_8130(clk,rst,matrix_A[8130],matrix_B[130],mul_res1[8130]);
multi_7x28 multi_7x28_mod_8131(clk,rst,matrix_A[8131],matrix_B[131],mul_res1[8131]);
multi_7x28 multi_7x28_mod_8132(clk,rst,matrix_A[8132],matrix_B[132],mul_res1[8132]);
multi_7x28 multi_7x28_mod_8133(clk,rst,matrix_A[8133],matrix_B[133],mul_res1[8133]);
multi_7x28 multi_7x28_mod_8134(clk,rst,matrix_A[8134],matrix_B[134],mul_res1[8134]);
multi_7x28 multi_7x28_mod_8135(clk,rst,matrix_A[8135],matrix_B[135],mul_res1[8135]);
multi_7x28 multi_7x28_mod_8136(clk,rst,matrix_A[8136],matrix_B[136],mul_res1[8136]);
multi_7x28 multi_7x28_mod_8137(clk,rst,matrix_A[8137],matrix_B[137],mul_res1[8137]);
multi_7x28 multi_7x28_mod_8138(clk,rst,matrix_A[8138],matrix_B[138],mul_res1[8138]);
multi_7x28 multi_7x28_mod_8139(clk,rst,matrix_A[8139],matrix_B[139],mul_res1[8139]);
multi_7x28 multi_7x28_mod_8140(clk,rst,matrix_A[8140],matrix_B[140],mul_res1[8140]);
multi_7x28 multi_7x28_mod_8141(clk,rst,matrix_A[8141],matrix_B[141],mul_res1[8141]);
multi_7x28 multi_7x28_mod_8142(clk,rst,matrix_A[8142],matrix_B[142],mul_res1[8142]);
multi_7x28 multi_7x28_mod_8143(clk,rst,matrix_A[8143],matrix_B[143],mul_res1[8143]);
multi_7x28 multi_7x28_mod_8144(clk,rst,matrix_A[8144],matrix_B[144],mul_res1[8144]);
multi_7x28 multi_7x28_mod_8145(clk,rst,matrix_A[8145],matrix_B[145],mul_res1[8145]);
multi_7x28 multi_7x28_mod_8146(clk,rst,matrix_A[8146],matrix_B[146],mul_res1[8146]);
multi_7x28 multi_7x28_mod_8147(clk,rst,matrix_A[8147],matrix_B[147],mul_res1[8147]);
multi_7x28 multi_7x28_mod_8148(clk,rst,matrix_A[8148],matrix_B[148],mul_res1[8148]);
multi_7x28 multi_7x28_mod_8149(clk,rst,matrix_A[8149],matrix_B[149],mul_res1[8149]);
multi_7x28 multi_7x28_mod_8150(clk,rst,matrix_A[8150],matrix_B[150],mul_res1[8150]);
multi_7x28 multi_7x28_mod_8151(clk,rst,matrix_A[8151],matrix_B[151],mul_res1[8151]);
multi_7x28 multi_7x28_mod_8152(clk,rst,matrix_A[8152],matrix_B[152],mul_res1[8152]);
multi_7x28 multi_7x28_mod_8153(clk,rst,matrix_A[8153],matrix_B[153],mul_res1[8153]);
multi_7x28 multi_7x28_mod_8154(clk,rst,matrix_A[8154],matrix_B[154],mul_res1[8154]);
multi_7x28 multi_7x28_mod_8155(clk,rst,matrix_A[8155],matrix_B[155],mul_res1[8155]);
multi_7x28 multi_7x28_mod_8156(clk,rst,matrix_A[8156],matrix_B[156],mul_res1[8156]);
multi_7x28 multi_7x28_mod_8157(clk,rst,matrix_A[8157],matrix_B[157],mul_res1[8157]);
multi_7x28 multi_7x28_mod_8158(clk,rst,matrix_A[8158],matrix_B[158],mul_res1[8158]);
multi_7x28 multi_7x28_mod_8159(clk,rst,matrix_A[8159],matrix_B[159],mul_res1[8159]);
multi_7x28 multi_7x28_mod_8160(clk,rst,matrix_A[8160],matrix_B[160],mul_res1[8160]);
multi_7x28 multi_7x28_mod_8161(clk,rst,matrix_A[8161],matrix_B[161],mul_res1[8161]);
multi_7x28 multi_7x28_mod_8162(clk,rst,matrix_A[8162],matrix_B[162],mul_res1[8162]);
multi_7x28 multi_7x28_mod_8163(clk,rst,matrix_A[8163],matrix_B[163],mul_res1[8163]);
multi_7x28 multi_7x28_mod_8164(clk,rst,matrix_A[8164],matrix_B[164],mul_res1[8164]);
multi_7x28 multi_7x28_mod_8165(clk,rst,matrix_A[8165],matrix_B[165],mul_res1[8165]);
multi_7x28 multi_7x28_mod_8166(clk,rst,matrix_A[8166],matrix_B[166],mul_res1[8166]);
multi_7x28 multi_7x28_mod_8167(clk,rst,matrix_A[8167],matrix_B[167],mul_res1[8167]);
multi_7x28 multi_7x28_mod_8168(clk,rst,matrix_A[8168],matrix_B[168],mul_res1[8168]);
multi_7x28 multi_7x28_mod_8169(clk,rst,matrix_A[8169],matrix_B[169],mul_res1[8169]);
multi_7x28 multi_7x28_mod_8170(clk,rst,matrix_A[8170],matrix_B[170],mul_res1[8170]);
multi_7x28 multi_7x28_mod_8171(clk,rst,matrix_A[8171],matrix_B[171],mul_res1[8171]);
multi_7x28 multi_7x28_mod_8172(clk,rst,matrix_A[8172],matrix_B[172],mul_res1[8172]);
multi_7x28 multi_7x28_mod_8173(clk,rst,matrix_A[8173],matrix_B[173],mul_res1[8173]);
multi_7x28 multi_7x28_mod_8174(clk,rst,matrix_A[8174],matrix_B[174],mul_res1[8174]);
multi_7x28 multi_7x28_mod_8175(clk,rst,matrix_A[8175],matrix_B[175],mul_res1[8175]);
multi_7x28 multi_7x28_mod_8176(clk,rst,matrix_A[8176],matrix_B[176],mul_res1[8176]);
multi_7x28 multi_7x28_mod_8177(clk,rst,matrix_A[8177],matrix_B[177],mul_res1[8177]);
multi_7x28 multi_7x28_mod_8178(clk,rst,matrix_A[8178],matrix_B[178],mul_res1[8178]);
multi_7x28 multi_7x28_mod_8179(clk,rst,matrix_A[8179],matrix_B[179],mul_res1[8179]);
multi_7x28 multi_7x28_mod_8180(clk,rst,matrix_A[8180],matrix_B[180],mul_res1[8180]);
multi_7x28 multi_7x28_mod_8181(clk,rst,matrix_A[8181],matrix_B[181],mul_res1[8181]);
multi_7x28 multi_7x28_mod_8182(clk,rst,matrix_A[8182],matrix_B[182],mul_res1[8182]);
multi_7x28 multi_7x28_mod_8183(clk,rst,matrix_A[8183],matrix_B[183],mul_res1[8183]);
multi_7x28 multi_7x28_mod_8184(clk,rst,matrix_A[8184],matrix_B[184],mul_res1[8184]);
multi_7x28 multi_7x28_mod_8185(clk,rst,matrix_A[8185],matrix_B[185],mul_res1[8185]);
multi_7x28 multi_7x28_mod_8186(clk,rst,matrix_A[8186],matrix_B[186],mul_res1[8186]);
multi_7x28 multi_7x28_mod_8187(clk,rst,matrix_A[8187],matrix_B[187],mul_res1[8187]);
multi_7x28 multi_7x28_mod_8188(clk,rst,matrix_A[8188],matrix_B[188],mul_res1[8188]);
multi_7x28 multi_7x28_mod_8189(clk,rst,matrix_A[8189],matrix_B[189],mul_res1[8189]);
multi_7x28 multi_7x28_mod_8190(clk,rst,matrix_A[8190],matrix_B[190],mul_res1[8190]);
multi_7x28 multi_7x28_mod_8191(clk,rst,matrix_A[8191],matrix_B[191],mul_res1[8191]);
multi_7x28 multi_7x28_mod_8192(clk,rst,matrix_A[8192],matrix_B[192],mul_res1[8192]);
multi_7x28 multi_7x28_mod_8193(clk,rst,matrix_A[8193],matrix_B[193],mul_res1[8193]);
multi_7x28 multi_7x28_mod_8194(clk,rst,matrix_A[8194],matrix_B[194],mul_res1[8194]);
multi_7x28 multi_7x28_mod_8195(clk,rst,matrix_A[8195],matrix_B[195],mul_res1[8195]);
multi_7x28 multi_7x28_mod_8196(clk,rst,matrix_A[8196],matrix_B[196],mul_res1[8196]);
multi_7x28 multi_7x28_mod_8197(clk,rst,matrix_A[8197],matrix_B[197],mul_res1[8197]);
multi_7x28 multi_7x28_mod_8198(clk,rst,matrix_A[8198],matrix_B[198],mul_res1[8198]);
multi_7x28 multi_7x28_mod_8199(clk,rst,matrix_A[8199],matrix_B[199],mul_res1[8199]);
multi_7x28 multi_7x28_mod_8200(clk,rst,matrix_A[8200],matrix_B[0],mul_res1[8200]);
multi_7x28 multi_7x28_mod_8201(clk,rst,matrix_A[8201],matrix_B[1],mul_res1[8201]);
multi_7x28 multi_7x28_mod_8202(clk,rst,matrix_A[8202],matrix_B[2],mul_res1[8202]);
multi_7x28 multi_7x28_mod_8203(clk,rst,matrix_A[8203],matrix_B[3],mul_res1[8203]);
multi_7x28 multi_7x28_mod_8204(clk,rst,matrix_A[8204],matrix_B[4],mul_res1[8204]);
multi_7x28 multi_7x28_mod_8205(clk,rst,matrix_A[8205],matrix_B[5],mul_res1[8205]);
multi_7x28 multi_7x28_mod_8206(clk,rst,matrix_A[8206],matrix_B[6],mul_res1[8206]);
multi_7x28 multi_7x28_mod_8207(clk,rst,matrix_A[8207],matrix_B[7],mul_res1[8207]);
multi_7x28 multi_7x28_mod_8208(clk,rst,matrix_A[8208],matrix_B[8],mul_res1[8208]);
multi_7x28 multi_7x28_mod_8209(clk,rst,matrix_A[8209],matrix_B[9],mul_res1[8209]);
multi_7x28 multi_7x28_mod_8210(clk,rst,matrix_A[8210],matrix_B[10],mul_res1[8210]);
multi_7x28 multi_7x28_mod_8211(clk,rst,matrix_A[8211],matrix_B[11],mul_res1[8211]);
multi_7x28 multi_7x28_mod_8212(clk,rst,matrix_A[8212],matrix_B[12],mul_res1[8212]);
multi_7x28 multi_7x28_mod_8213(clk,rst,matrix_A[8213],matrix_B[13],mul_res1[8213]);
multi_7x28 multi_7x28_mod_8214(clk,rst,matrix_A[8214],matrix_B[14],mul_res1[8214]);
multi_7x28 multi_7x28_mod_8215(clk,rst,matrix_A[8215],matrix_B[15],mul_res1[8215]);
multi_7x28 multi_7x28_mod_8216(clk,rst,matrix_A[8216],matrix_B[16],mul_res1[8216]);
multi_7x28 multi_7x28_mod_8217(clk,rst,matrix_A[8217],matrix_B[17],mul_res1[8217]);
multi_7x28 multi_7x28_mod_8218(clk,rst,matrix_A[8218],matrix_B[18],mul_res1[8218]);
multi_7x28 multi_7x28_mod_8219(clk,rst,matrix_A[8219],matrix_B[19],mul_res1[8219]);
multi_7x28 multi_7x28_mod_8220(clk,rst,matrix_A[8220],matrix_B[20],mul_res1[8220]);
multi_7x28 multi_7x28_mod_8221(clk,rst,matrix_A[8221],matrix_B[21],mul_res1[8221]);
multi_7x28 multi_7x28_mod_8222(clk,rst,matrix_A[8222],matrix_B[22],mul_res1[8222]);
multi_7x28 multi_7x28_mod_8223(clk,rst,matrix_A[8223],matrix_B[23],mul_res1[8223]);
multi_7x28 multi_7x28_mod_8224(clk,rst,matrix_A[8224],matrix_B[24],mul_res1[8224]);
multi_7x28 multi_7x28_mod_8225(clk,rst,matrix_A[8225],matrix_B[25],mul_res1[8225]);
multi_7x28 multi_7x28_mod_8226(clk,rst,matrix_A[8226],matrix_B[26],mul_res1[8226]);
multi_7x28 multi_7x28_mod_8227(clk,rst,matrix_A[8227],matrix_B[27],mul_res1[8227]);
multi_7x28 multi_7x28_mod_8228(clk,rst,matrix_A[8228],matrix_B[28],mul_res1[8228]);
multi_7x28 multi_7x28_mod_8229(clk,rst,matrix_A[8229],matrix_B[29],mul_res1[8229]);
multi_7x28 multi_7x28_mod_8230(clk,rst,matrix_A[8230],matrix_B[30],mul_res1[8230]);
multi_7x28 multi_7x28_mod_8231(clk,rst,matrix_A[8231],matrix_B[31],mul_res1[8231]);
multi_7x28 multi_7x28_mod_8232(clk,rst,matrix_A[8232],matrix_B[32],mul_res1[8232]);
multi_7x28 multi_7x28_mod_8233(clk,rst,matrix_A[8233],matrix_B[33],mul_res1[8233]);
multi_7x28 multi_7x28_mod_8234(clk,rst,matrix_A[8234],matrix_B[34],mul_res1[8234]);
multi_7x28 multi_7x28_mod_8235(clk,rst,matrix_A[8235],matrix_B[35],mul_res1[8235]);
multi_7x28 multi_7x28_mod_8236(clk,rst,matrix_A[8236],matrix_B[36],mul_res1[8236]);
multi_7x28 multi_7x28_mod_8237(clk,rst,matrix_A[8237],matrix_B[37],mul_res1[8237]);
multi_7x28 multi_7x28_mod_8238(clk,rst,matrix_A[8238],matrix_B[38],mul_res1[8238]);
multi_7x28 multi_7x28_mod_8239(clk,rst,matrix_A[8239],matrix_B[39],mul_res1[8239]);
multi_7x28 multi_7x28_mod_8240(clk,rst,matrix_A[8240],matrix_B[40],mul_res1[8240]);
multi_7x28 multi_7x28_mod_8241(clk,rst,matrix_A[8241],matrix_B[41],mul_res1[8241]);
multi_7x28 multi_7x28_mod_8242(clk,rst,matrix_A[8242],matrix_B[42],mul_res1[8242]);
multi_7x28 multi_7x28_mod_8243(clk,rst,matrix_A[8243],matrix_B[43],mul_res1[8243]);
multi_7x28 multi_7x28_mod_8244(clk,rst,matrix_A[8244],matrix_B[44],mul_res1[8244]);
multi_7x28 multi_7x28_mod_8245(clk,rst,matrix_A[8245],matrix_B[45],mul_res1[8245]);
multi_7x28 multi_7x28_mod_8246(clk,rst,matrix_A[8246],matrix_B[46],mul_res1[8246]);
multi_7x28 multi_7x28_mod_8247(clk,rst,matrix_A[8247],matrix_B[47],mul_res1[8247]);
multi_7x28 multi_7x28_mod_8248(clk,rst,matrix_A[8248],matrix_B[48],mul_res1[8248]);
multi_7x28 multi_7x28_mod_8249(clk,rst,matrix_A[8249],matrix_B[49],mul_res1[8249]);
multi_7x28 multi_7x28_mod_8250(clk,rst,matrix_A[8250],matrix_B[50],mul_res1[8250]);
multi_7x28 multi_7x28_mod_8251(clk,rst,matrix_A[8251],matrix_B[51],mul_res1[8251]);
multi_7x28 multi_7x28_mod_8252(clk,rst,matrix_A[8252],matrix_B[52],mul_res1[8252]);
multi_7x28 multi_7x28_mod_8253(clk,rst,matrix_A[8253],matrix_B[53],mul_res1[8253]);
multi_7x28 multi_7x28_mod_8254(clk,rst,matrix_A[8254],matrix_B[54],mul_res1[8254]);
multi_7x28 multi_7x28_mod_8255(clk,rst,matrix_A[8255],matrix_B[55],mul_res1[8255]);
multi_7x28 multi_7x28_mod_8256(clk,rst,matrix_A[8256],matrix_B[56],mul_res1[8256]);
multi_7x28 multi_7x28_mod_8257(clk,rst,matrix_A[8257],matrix_B[57],mul_res1[8257]);
multi_7x28 multi_7x28_mod_8258(clk,rst,matrix_A[8258],matrix_B[58],mul_res1[8258]);
multi_7x28 multi_7x28_mod_8259(clk,rst,matrix_A[8259],matrix_B[59],mul_res1[8259]);
multi_7x28 multi_7x28_mod_8260(clk,rst,matrix_A[8260],matrix_B[60],mul_res1[8260]);
multi_7x28 multi_7x28_mod_8261(clk,rst,matrix_A[8261],matrix_B[61],mul_res1[8261]);
multi_7x28 multi_7x28_mod_8262(clk,rst,matrix_A[8262],matrix_B[62],mul_res1[8262]);
multi_7x28 multi_7x28_mod_8263(clk,rst,matrix_A[8263],matrix_B[63],mul_res1[8263]);
multi_7x28 multi_7x28_mod_8264(clk,rst,matrix_A[8264],matrix_B[64],mul_res1[8264]);
multi_7x28 multi_7x28_mod_8265(clk,rst,matrix_A[8265],matrix_B[65],mul_res1[8265]);
multi_7x28 multi_7x28_mod_8266(clk,rst,matrix_A[8266],matrix_B[66],mul_res1[8266]);
multi_7x28 multi_7x28_mod_8267(clk,rst,matrix_A[8267],matrix_B[67],mul_res1[8267]);
multi_7x28 multi_7x28_mod_8268(clk,rst,matrix_A[8268],matrix_B[68],mul_res1[8268]);
multi_7x28 multi_7x28_mod_8269(clk,rst,matrix_A[8269],matrix_B[69],mul_res1[8269]);
multi_7x28 multi_7x28_mod_8270(clk,rst,matrix_A[8270],matrix_B[70],mul_res1[8270]);
multi_7x28 multi_7x28_mod_8271(clk,rst,matrix_A[8271],matrix_B[71],mul_res1[8271]);
multi_7x28 multi_7x28_mod_8272(clk,rst,matrix_A[8272],matrix_B[72],mul_res1[8272]);
multi_7x28 multi_7x28_mod_8273(clk,rst,matrix_A[8273],matrix_B[73],mul_res1[8273]);
multi_7x28 multi_7x28_mod_8274(clk,rst,matrix_A[8274],matrix_B[74],mul_res1[8274]);
multi_7x28 multi_7x28_mod_8275(clk,rst,matrix_A[8275],matrix_B[75],mul_res1[8275]);
multi_7x28 multi_7x28_mod_8276(clk,rst,matrix_A[8276],matrix_B[76],mul_res1[8276]);
multi_7x28 multi_7x28_mod_8277(clk,rst,matrix_A[8277],matrix_B[77],mul_res1[8277]);
multi_7x28 multi_7x28_mod_8278(clk,rst,matrix_A[8278],matrix_B[78],mul_res1[8278]);
multi_7x28 multi_7x28_mod_8279(clk,rst,matrix_A[8279],matrix_B[79],mul_res1[8279]);
multi_7x28 multi_7x28_mod_8280(clk,rst,matrix_A[8280],matrix_B[80],mul_res1[8280]);
multi_7x28 multi_7x28_mod_8281(clk,rst,matrix_A[8281],matrix_B[81],mul_res1[8281]);
multi_7x28 multi_7x28_mod_8282(clk,rst,matrix_A[8282],matrix_B[82],mul_res1[8282]);
multi_7x28 multi_7x28_mod_8283(clk,rst,matrix_A[8283],matrix_B[83],mul_res1[8283]);
multi_7x28 multi_7x28_mod_8284(clk,rst,matrix_A[8284],matrix_B[84],mul_res1[8284]);
multi_7x28 multi_7x28_mod_8285(clk,rst,matrix_A[8285],matrix_B[85],mul_res1[8285]);
multi_7x28 multi_7x28_mod_8286(clk,rst,matrix_A[8286],matrix_B[86],mul_res1[8286]);
multi_7x28 multi_7x28_mod_8287(clk,rst,matrix_A[8287],matrix_B[87],mul_res1[8287]);
multi_7x28 multi_7x28_mod_8288(clk,rst,matrix_A[8288],matrix_B[88],mul_res1[8288]);
multi_7x28 multi_7x28_mod_8289(clk,rst,matrix_A[8289],matrix_B[89],mul_res1[8289]);
multi_7x28 multi_7x28_mod_8290(clk,rst,matrix_A[8290],matrix_B[90],mul_res1[8290]);
multi_7x28 multi_7x28_mod_8291(clk,rst,matrix_A[8291],matrix_B[91],mul_res1[8291]);
multi_7x28 multi_7x28_mod_8292(clk,rst,matrix_A[8292],matrix_B[92],mul_res1[8292]);
multi_7x28 multi_7x28_mod_8293(clk,rst,matrix_A[8293],matrix_B[93],mul_res1[8293]);
multi_7x28 multi_7x28_mod_8294(clk,rst,matrix_A[8294],matrix_B[94],mul_res1[8294]);
multi_7x28 multi_7x28_mod_8295(clk,rst,matrix_A[8295],matrix_B[95],mul_res1[8295]);
multi_7x28 multi_7x28_mod_8296(clk,rst,matrix_A[8296],matrix_B[96],mul_res1[8296]);
multi_7x28 multi_7x28_mod_8297(clk,rst,matrix_A[8297],matrix_B[97],mul_res1[8297]);
multi_7x28 multi_7x28_mod_8298(clk,rst,matrix_A[8298],matrix_B[98],mul_res1[8298]);
multi_7x28 multi_7x28_mod_8299(clk,rst,matrix_A[8299],matrix_B[99],mul_res1[8299]);
multi_7x28 multi_7x28_mod_8300(clk,rst,matrix_A[8300],matrix_B[100],mul_res1[8300]);
multi_7x28 multi_7x28_mod_8301(clk,rst,matrix_A[8301],matrix_B[101],mul_res1[8301]);
multi_7x28 multi_7x28_mod_8302(clk,rst,matrix_A[8302],matrix_B[102],mul_res1[8302]);
multi_7x28 multi_7x28_mod_8303(clk,rst,matrix_A[8303],matrix_B[103],mul_res1[8303]);
multi_7x28 multi_7x28_mod_8304(clk,rst,matrix_A[8304],matrix_B[104],mul_res1[8304]);
multi_7x28 multi_7x28_mod_8305(clk,rst,matrix_A[8305],matrix_B[105],mul_res1[8305]);
multi_7x28 multi_7x28_mod_8306(clk,rst,matrix_A[8306],matrix_B[106],mul_res1[8306]);
multi_7x28 multi_7x28_mod_8307(clk,rst,matrix_A[8307],matrix_B[107],mul_res1[8307]);
multi_7x28 multi_7x28_mod_8308(clk,rst,matrix_A[8308],matrix_B[108],mul_res1[8308]);
multi_7x28 multi_7x28_mod_8309(clk,rst,matrix_A[8309],matrix_B[109],mul_res1[8309]);
multi_7x28 multi_7x28_mod_8310(clk,rst,matrix_A[8310],matrix_B[110],mul_res1[8310]);
multi_7x28 multi_7x28_mod_8311(clk,rst,matrix_A[8311],matrix_B[111],mul_res1[8311]);
multi_7x28 multi_7x28_mod_8312(clk,rst,matrix_A[8312],matrix_B[112],mul_res1[8312]);
multi_7x28 multi_7x28_mod_8313(clk,rst,matrix_A[8313],matrix_B[113],mul_res1[8313]);
multi_7x28 multi_7x28_mod_8314(clk,rst,matrix_A[8314],matrix_B[114],mul_res1[8314]);
multi_7x28 multi_7x28_mod_8315(clk,rst,matrix_A[8315],matrix_B[115],mul_res1[8315]);
multi_7x28 multi_7x28_mod_8316(clk,rst,matrix_A[8316],matrix_B[116],mul_res1[8316]);
multi_7x28 multi_7x28_mod_8317(clk,rst,matrix_A[8317],matrix_B[117],mul_res1[8317]);
multi_7x28 multi_7x28_mod_8318(clk,rst,matrix_A[8318],matrix_B[118],mul_res1[8318]);
multi_7x28 multi_7x28_mod_8319(clk,rst,matrix_A[8319],matrix_B[119],mul_res1[8319]);
multi_7x28 multi_7x28_mod_8320(clk,rst,matrix_A[8320],matrix_B[120],mul_res1[8320]);
multi_7x28 multi_7x28_mod_8321(clk,rst,matrix_A[8321],matrix_B[121],mul_res1[8321]);
multi_7x28 multi_7x28_mod_8322(clk,rst,matrix_A[8322],matrix_B[122],mul_res1[8322]);
multi_7x28 multi_7x28_mod_8323(clk,rst,matrix_A[8323],matrix_B[123],mul_res1[8323]);
multi_7x28 multi_7x28_mod_8324(clk,rst,matrix_A[8324],matrix_B[124],mul_res1[8324]);
multi_7x28 multi_7x28_mod_8325(clk,rst,matrix_A[8325],matrix_B[125],mul_res1[8325]);
multi_7x28 multi_7x28_mod_8326(clk,rst,matrix_A[8326],matrix_B[126],mul_res1[8326]);
multi_7x28 multi_7x28_mod_8327(clk,rst,matrix_A[8327],matrix_B[127],mul_res1[8327]);
multi_7x28 multi_7x28_mod_8328(clk,rst,matrix_A[8328],matrix_B[128],mul_res1[8328]);
multi_7x28 multi_7x28_mod_8329(clk,rst,matrix_A[8329],matrix_B[129],mul_res1[8329]);
multi_7x28 multi_7x28_mod_8330(clk,rst,matrix_A[8330],matrix_B[130],mul_res1[8330]);
multi_7x28 multi_7x28_mod_8331(clk,rst,matrix_A[8331],matrix_B[131],mul_res1[8331]);
multi_7x28 multi_7x28_mod_8332(clk,rst,matrix_A[8332],matrix_B[132],mul_res1[8332]);
multi_7x28 multi_7x28_mod_8333(clk,rst,matrix_A[8333],matrix_B[133],mul_res1[8333]);
multi_7x28 multi_7x28_mod_8334(clk,rst,matrix_A[8334],matrix_B[134],mul_res1[8334]);
multi_7x28 multi_7x28_mod_8335(clk,rst,matrix_A[8335],matrix_B[135],mul_res1[8335]);
multi_7x28 multi_7x28_mod_8336(clk,rst,matrix_A[8336],matrix_B[136],mul_res1[8336]);
multi_7x28 multi_7x28_mod_8337(clk,rst,matrix_A[8337],matrix_B[137],mul_res1[8337]);
multi_7x28 multi_7x28_mod_8338(clk,rst,matrix_A[8338],matrix_B[138],mul_res1[8338]);
multi_7x28 multi_7x28_mod_8339(clk,rst,matrix_A[8339],matrix_B[139],mul_res1[8339]);
multi_7x28 multi_7x28_mod_8340(clk,rst,matrix_A[8340],matrix_B[140],mul_res1[8340]);
multi_7x28 multi_7x28_mod_8341(clk,rst,matrix_A[8341],matrix_B[141],mul_res1[8341]);
multi_7x28 multi_7x28_mod_8342(clk,rst,matrix_A[8342],matrix_B[142],mul_res1[8342]);
multi_7x28 multi_7x28_mod_8343(clk,rst,matrix_A[8343],matrix_B[143],mul_res1[8343]);
multi_7x28 multi_7x28_mod_8344(clk,rst,matrix_A[8344],matrix_B[144],mul_res1[8344]);
multi_7x28 multi_7x28_mod_8345(clk,rst,matrix_A[8345],matrix_B[145],mul_res1[8345]);
multi_7x28 multi_7x28_mod_8346(clk,rst,matrix_A[8346],matrix_B[146],mul_res1[8346]);
multi_7x28 multi_7x28_mod_8347(clk,rst,matrix_A[8347],matrix_B[147],mul_res1[8347]);
multi_7x28 multi_7x28_mod_8348(clk,rst,matrix_A[8348],matrix_B[148],mul_res1[8348]);
multi_7x28 multi_7x28_mod_8349(clk,rst,matrix_A[8349],matrix_B[149],mul_res1[8349]);
multi_7x28 multi_7x28_mod_8350(clk,rst,matrix_A[8350],matrix_B[150],mul_res1[8350]);
multi_7x28 multi_7x28_mod_8351(clk,rst,matrix_A[8351],matrix_B[151],mul_res1[8351]);
multi_7x28 multi_7x28_mod_8352(clk,rst,matrix_A[8352],matrix_B[152],mul_res1[8352]);
multi_7x28 multi_7x28_mod_8353(clk,rst,matrix_A[8353],matrix_B[153],mul_res1[8353]);
multi_7x28 multi_7x28_mod_8354(clk,rst,matrix_A[8354],matrix_B[154],mul_res1[8354]);
multi_7x28 multi_7x28_mod_8355(clk,rst,matrix_A[8355],matrix_B[155],mul_res1[8355]);
multi_7x28 multi_7x28_mod_8356(clk,rst,matrix_A[8356],matrix_B[156],mul_res1[8356]);
multi_7x28 multi_7x28_mod_8357(clk,rst,matrix_A[8357],matrix_B[157],mul_res1[8357]);
multi_7x28 multi_7x28_mod_8358(clk,rst,matrix_A[8358],matrix_B[158],mul_res1[8358]);
multi_7x28 multi_7x28_mod_8359(clk,rst,matrix_A[8359],matrix_B[159],mul_res1[8359]);
multi_7x28 multi_7x28_mod_8360(clk,rst,matrix_A[8360],matrix_B[160],mul_res1[8360]);
multi_7x28 multi_7x28_mod_8361(clk,rst,matrix_A[8361],matrix_B[161],mul_res1[8361]);
multi_7x28 multi_7x28_mod_8362(clk,rst,matrix_A[8362],matrix_B[162],mul_res1[8362]);
multi_7x28 multi_7x28_mod_8363(clk,rst,matrix_A[8363],matrix_B[163],mul_res1[8363]);
multi_7x28 multi_7x28_mod_8364(clk,rst,matrix_A[8364],matrix_B[164],mul_res1[8364]);
multi_7x28 multi_7x28_mod_8365(clk,rst,matrix_A[8365],matrix_B[165],mul_res1[8365]);
multi_7x28 multi_7x28_mod_8366(clk,rst,matrix_A[8366],matrix_B[166],mul_res1[8366]);
multi_7x28 multi_7x28_mod_8367(clk,rst,matrix_A[8367],matrix_B[167],mul_res1[8367]);
multi_7x28 multi_7x28_mod_8368(clk,rst,matrix_A[8368],matrix_B[168],mul_res1[8368]);
multi_7x28 multi_7x28_mod_8369(clk,rst,matrix_A[8369],matrix_B[169],mul_res1[8369]);
multi_7x28 multi_7x28_mod_8370(clk,rst,matrix_A[8370],matrix_B[170],mul_res1[8370]);
multi_7x28 multi_7x28_mod_8371(clk,rst,matrix_A[8371],matrix_B[171],mul_res1[8371]);
multi_7x28 multi_7x28_mod_8372(clk,rst,matrix_A[8372],matrix_B[172],mul_res1[8372]);
multi_7x28 multi_7x28_mod_8373(clk,rst,matrix_A[8373],matrix_B[173],mul_res1[8373]);
multi_7x28 multi_7x28_mod_8374(clk,rst,matrix_A[8374],matrix_B[174],mul_res1[8374]);
multi_7x28 multi_7x28_mod_8375(clk,rst,matrix_A[8375],matrix_B[175],mul_res1[8375]);
multi_7x28 multi_7x28_mod_8376(clk,rst,matrix_A[8376],matrix_B[176],mul_res1[8376]);
multi_7x28 multi_7x28_mod_8377(clk,rst,matrix_A[8377],matrix_B[177],mul_res1[8377]);
multi_7x28 multi_7x28_mod_8378(clk,rst,matrix_A[8378],matrix_B[178],mul_res1[8378]);
multi_7x28 multi_7x28_mod_8379(clk,rst,matrix_A[8379],matrix_B[179],mul_res1[8379]);
multi_7x28 multi_7x28_mod_8380(clk,rst,matrix_A[8380],matrix_B[180],mul_res1[8380]);
multi_7x28 multi_7x28_mod_8381(clk,rst,matrix_A[8381],matrix_B[181],mul_res1[8381]);
multi_7x28 multi_7x28_mod_8382(clk,rst,matrix_A[8382],matrix_B[182],mul_res1[8382]);
multi_7x28 multi_7x28_mod_8383(clk,rst,matrix_A[8383],matrix_B[183],mul_res1[8383]);
multi_7x28 multi_7x28_mod_8384(clk,rst,matrix_A[8384],matrix_B[184],mul_res1[8384]);
multi_7x28 multi_7x28_mod_8385(clk,rst,matrix_A[8385],matrix_B[185],mul_res1[8385]);
multi_7x28 multi_7x28_mod_8386(clk,rst,matrix_A[8386],matrix_B[186],mul_res1[8386]);
multi_7x28 multi_7x28_mod_8387(clk,rst,matrix_A[8387],matrix_B[187],mul_res1[8387]);
multi_7x28 multi_7x28_mod_8388(clk,rst,matrix_A[8388],matrix_B[188],mul_res1[8388]);
multi_7x28 multi_7x28_mod_8389(clk,rst,matrix_A[8389],matrix_B[189],mul_res1[8389]);
multi_7x28 multi_7x28_mod_8390(clk,rst,matrix_A[8390],matrix_B[190],mul_res1[8390]);
multi_7x28 multi_7x28_mod_8391(clk,rst,matrix_A[8391],matrix_B[191],mul_res1[8391]);
multi_7x28 multi_7x28_mod_8392(clk,rst,matrix_A[8392],matrix_B[192],mul_res1[8392]);
multi_7x28 multi_7x28_mod_8393(clk,rst,matrix_A[8393],matrix_B[193],mul_res1[8393]);
multi_7x28 multi_7x28_mod_8394(clk,rst,matrix_A[8394],matrix_B[194],mul_res1[8394]);
multi_7x28 multi_7x28_mod_8395(clk,rst,matrix_A[8395],matrix_B[195],mul_res1[8395]);
multi_7x28 multi_7x28_mod_8396(clk,rst,matrix_A[8396],matrix_B[196],mul_res1[8396]);
multi_7x28 multi_7x28_mod_8397(clk,rst,matrix_A[8397],matrix_B[197],mul_res1[8397]);
multi_7x28 multi_7x28_mod_8398(clk,rst,matrix_A[8398],matrix_B[198],mul_res1[8398]);
multi_7x28 multi_7x28_mod_8399(clk,rst,matrix_A[8399],matrix_B[199],mul_res1[8399]);
multi_7x28 multi_7x28_mod_8400(clk,rst,matrix_A[8400],matrix_B[0],mul_res1[8400]);
multi_7x28 multi_7x28_mod_8401(clk,rst,matrix_A[8401],matrix_B[1],mul_res1[8401]);
multi_7x28 multi_7x28_mod_8402(clk,rst,matrix_A[8402],matrix_B[2],mul_res1[8402]);
multi_7x28 multi_7x28_mod_8403(clk,rst,matrix_A[8403],matrix_B[3],mul_res1[8403]);
multi_7x28 multi_7x28_mod_8404(clk,rst,matrix_A[8404],matrix_B[4],mul_res1[8404]);
multi_7x28 multi_7x28_mod_8405(clk,rst,matrix_A[8405],matrix_B[5],mul_res1[8405]);
multi_7x28 multi_7x28_mod_8406(clk,rst,matrix_A[8406],matrix_B[6],mul_res1[8406]);
multi_7x28 multi_7x28_mod_8407(clk,rst,matrix_A[8407],matrix_B[7],mul_res1[8407]);
multi_7x28 multi_7x28_mod_8408(clk,rst,matrix_A[8408],matrix_B[8],mul_res1[8408]);
multi_7x28 multi_7x28_mod_8409(clk,rst,matrix_A[8409],matrix_B[9],mul_res1[8409]);
multi_7x28 multi_7x28_mod_8410(clk,rst,matrix_A[8410],matrix_B[10],mul_res1[8410]);
multi_7x28 multi_7x28_mod_8411(clk,rst,matrix_A[8411],matrix_B[11],mul_res1[8411]);
multi_7x28 multi_7x28_mod_8412(clk,rst,matrix_A[8412],matrix_B[12],mul_res1[8412]);
multi_7x28 multi_7x28_mod_8413(clk,rst,matrix_A[8413],matrix_B[13],mul_res1[8413]);
multi_7x28 multi_7x28_mod_8414(clk,rst,matrix_A[8414],matrix_B[14],mul_res1[8414]);
multi_7x28 multi_7x28_mod_8415(clk,rst,matrix_A[8415],matrix_B[15],mul_res1[8415]);
multi_7x28 multi_7x28_mod_8416(clk,rst,matrix_A[8416],matrix_B[16],mul_res1[8416]);
multi_7x28 multi_7x28_mod_8417(clk,rst,matrix_A[8417],matrix_B[17],mul_res1[8417]);
multi_7x28 multi_7x28_mod_8418(clk,rst,matrix_A[8418],matrix_B[18],mul_res1[8418]);
multi_7x28 multi_7x28_mod_8419(clk,rst,matrix_A[8419],matrix_B[19],mul_res1[8419]);
multi_7x28 multi_7x28_mod_8420(clk,rst,matrix_A[8420],matrix_B[20],mul_res1[8420]);
multi_7x28 multi_7x28_mod_8421(clk,rst,matrix_A[8421],matrix_B[21],mul_res1[8421]);
multi_7x28 multi_7x28_mod_8422(clk,rst,matrix_A[8422],matrix_B[22],mul_res1[8422]);
multi_7x28 multi_7x28_mod_8423(clk,rst,matrix_A[8423],matrix_B[23],mul_res1[8423]);
multi_7x28 multi_7x28_mod_8424(clk,rst,matrix_A[8424],matrix_B[24],mul_res1[8424]);
multi_7x28 multi_7x28_mod_8425(clk,rst,matrix_A[8425],matrix_B[25],mul_res1[8425]);
multi_7x28 multi_7x28_mod_8426(clk,rst,matrix_A[8426],matrix_B[26],mul_res1[8426]);
multi_7x28 multi_7x28_mod_8427(clk,rst,matrix_A[8427],matrix_B[27],mul_res1[8427]);
multi_7x28 multi_7x28_mod_8428(clk,rst,matrix_A[8428],matrix_B[28],mul_res1[8428]);
multi_7x28 multi_7x28_mod_8429(clk,rst,matrix_A[8429],matrix_B[29],mul_res1[8429]);
multi_7x28 multi_7x28_mod_8430(clk,rst,matrix_A[8430],matrix_B[30],mul_res1[8430]);
multi_7x28 multi_7x28_mod_8431(clk,rst,matrix_A[8431],matrix_B[31],mul_res1[8431]);
multi_7x28 multi_7x28_mod_8432(clk,rst,matrix_A[8432],matrix_B[32],mul_res1[8432]);
multi_7x28 multi_7x28_mod_8433(clk,rst,matrix_A[8433],matrix_B[33],mul_res1[8433]);
multi_7x28 multi_7x28_mod_8434(clk,rst,matrix_A[8434],matrix_B[34],mul_res1[8434]);
multi_7x28 multi_7x28_mod_8435(clk,rst,matrix_A[8435],matrix_B[35],mul_res1[8435]);
multi_7x28 multi_7x28_mod_8436(clk,rst,matrix_A[8436],matrix_B[36],mul_res1[8436]);
multi_7x28 multi_7x28_mod_8437(clk,rst,matrix_A[8437],matrix_B[37],mul_res1[8437]);
multi_7x28 multi_7x28_mod_8438(clk,rst,matrix_A[8438],matrix_B[38],mul_res1[8438]);
multi_7x28 multi_7x28_mod_8439(clk,rst,matrix_A[8439],matrix_B[39],mul_res1[8439]);
multi_7x28 multi_7x28_mod_8440(clk,rst,matrix_A[8440],matrix_B[40],mul_res1[8440]);
multi_7x28 multi_7x28_mod_8441(clk,rst,matrix_A[8441],matrix_B[41],mul_res1[8441]);
multi_7x28 multi_7x28_mod_8442(clk,rst,matrix_A[8442],matrix_B[42],mul_res1[8442]);
multi_7x28 multi_7x28_mod_8443(clk,rst,matrix_A[8443],matrix_B[43],mul_res1[8443]);
multi_7x28 multi_7x28_mod_8444(clk,rst,matrix_A[8444],matrix_B[44],mul_res1[8444]);
multi_7x28 multi_7x28_mod_8445(clk,rst,matrix_A[8445],matrix_B[45],mul_res1[8445]);
multi_7x28 multi_7x28_mod_8446(clk,rst,matrix_A[8446],matrix_B[46],mul_res1[8446]);
multi_7x28 multi_7x28_mod_8447(clk,rst,matrix_A[8447],matrix_B[47],mul_res1[8447]);
multi_7x28 multi_7x28_mod_8448(clk,rst,matrix_A[8448],matrix_B[48],mul_res1[8448]);
multi_7x28 multi_7x28_mod_8449(clk,rst,matrix_A[8449],matrix_B[49],mul_res1[8449]);
multi_7x28 multi_7x28_mod_8450(clk,rst,matrix_A[8450],matrix_B[50],mul_res1[8450]);
multi_7x28 multi_7x28_mod_8451(clk,rst,matrix_A[8451],matrix_B[51],mul_res1[8451]);
multi_7x28 multi_7x28_mod_8452(clk,rst,matrix_A[8452],matrix_B[52],mul_res1[8452]);
multi_7x28 multi_7x28_mod_8453(clk,rst,matrix_A[8453],matrix_B[53],mul_res1[8453]);
multi_7x28 multi_7x28_mod_8454(clk,rst,matrix_A[8454],matrix_B[54],mul_res1[8454]);
multi_7x28 multi_7x28_mod_8455(clk,rst,matrix_A[8455],matrix_B[55],mul_res1[8455]);
multi_7x28 multi_7x28_mod_8456(clk,rst,matrix_A[8456],matrix_B[56],mul_res1[8456]);
multi_7x28 multi_7x28_mod_8457(clk,rst,matrix_A[8457],matrix_B[57],mul_res1[8457]);
multi_7x28 multi_7x28_mod_8458(clk,rst,matrix_A[8458],matrix_B[58],mul_res1[8458]);
multi_7x28 multi_7x28_mod_8459(clk,rst,matrix_A[8459],matrix_B[59],mul_res1[8459]);
multi_7x28 multi_7x28_mod_8460(clk,rst,matrix_A[8460],matrix_B[60],mul_res1[8460]);
multi_7x28 multi_7x28_mod_8461(clk,rst,matrix_A[8461],matrix_B[61],mul_res1[8461]);
multi_7x28 multi_7x28_mod_8462(clk,rst,matrix_A[8462],matrix_B[62],mul_res1[8462]);
multi_7x28 multi_7x28_mod_8463(clk,rst,matrix_A[8463],matrix_B[63],mul_res1[8463]);
multi_7x28 multi_7x28_mod_8464(clk,rst,matrix_A[8464],matrix_B[64],mul_res1[8464]);
multi_7x28 multi_7x28_mod_8465(clk,rst,matrix_A[8465],matrix_B[65],mul_res1[8465]);
multi_7x28 multi_7x28_mod_8466(clk,rst,matrix_A[8466],matrix_B[66],mul_res1[8466]);
multi_7x28 multi_7x28_mod_8467(clk,rst,matrix_A[8467],matrix_B[67],mul_res1[8467]);
multi_7x28 multi_7x28_mod_8468(clk,rst,matrix_A[8468],matrix_B[68],mul_res1[8468]);
multi_7x28 multi_7x28_mod_8469(clk,rst,matrix_A[8469],matrix_B[69],mul_res1[8469]);
multi_7x28 multi_7x28_mod_8470(clk,rst,matrix_A[8470],matrix_B[70],mul_res1[8470]);
multi_7x28 multi_7x28_mod_8471(clk,rst,matrix_A[8471],matrix_B[71],mul_res1[8471]);
multi_7x28 multi_7x28_mod_8472(clk,rst,matrix_A[8472],matrix_B[72],mul_res1[8472]);
multi_7x28 multi_7x28_mod_8473(clk,rst,matrix_A[8473],matrix_B[73],mul_res1[8473]);
multi_7x28 multi_7x28_mod_8474(clk,rst,matrix_A[8474],matrix_B[74],mul_res1[8474]);
multi_7x28 multi_7x28_mod_8475(clk,rst,matrix_A[8475],matrix_B[75],mul_res1[8475]);
multi_7x28 multi_7x28_mod_8476(clk,rst,matrix_A[8476],matrix_B[76],mul_res1[8476]);
multi_7x28 multi_7x28_mod_8477(clk,rst,matrix_A[8477],matrix_B[77],mul_res1[8477]);
multi_7x28 multi_7x28_mod_8478(clk,rst,matrix_A[8478],matrix_B[78],mul_res1[8478]);
multi_7x28 multi_7x28_mod_8479(clk,rst,matrix_A[8479],matrix_B[79],mul_res1[8479]);
multi_7x28 multi_7x28_mod_8480(clk,rst,matrix_A[8480],matrix_B[80],mul_res1[8480]);
multi_7x28 multi_7x28_mod_8481(clk,rst,matrix_A[8481],matrix_B[81],mul_res1[8481]);
multi_7x28 multi_7x28_mod_8482(clk,rst,matrix_A[8482],matrix_B[82],mul_res1[8482]);
multi_7x28 multi_7x28_mod_8483(clk,rst,matrix_A[8483],matrix_B[83],mul_res1[8483]);
multi_7x28 multi_7x28_mod_8484(clk,rst,matrix_A[8484],matrix_B[84],mul_res1[8484]);
multi_7x28 multi_7x28_mod_8485(clk,rst,matrix_A[8485],matrix_B[85],mul_res1[8485]);
multi_7x28 multi_7x28_mod_8486(clk,rst,matrix_A[8486],matrix_B[86],mul_res1[8486]);
multi_7x28 multi_7x28_mod_8487(clk,rst,matrix_A[8487],matrix_B[87],mul_res1[8487]);
multi_7x28 multi_7x28_mod_8488(clk,rst,matrix_A[8488],matrix_B[88],mul_res1[8488]);
multi_7x28 multi_7x28_mod_8489(clk,rst,matrix_A[8489],matrix_B[89],mul_res1[8489]);
multi_7x28 multi_7x28_mod_8490(clk,rst,matrix_A[8490],matrix_B[90],mul_res1[8490]);
multi_7x28 multi_7x28_mod_8491(clk,rst,matrix_A[8491],matrix_B[91],mul_res1[8491]);
multi_7x28 multi_7x28_mod_8492(clk,rst,matrix_A[8492],matrix_B[92],mul_res1[8492]);
multi_7x28 multi_7x28_mod_8493(clk,rst,matrix_A[8493],matrix_B[93],mul_res1[8493]);
multi_7x28 multi_7x28_mod_8494(clk,rst,matrix_A[8494],matrix_B[94],mul_res1[8494]);
multi_7x28 multi_7x28_mod_8495(clk,rst,matrix_A[8495],matrix_B[95],mul_res1[8495]);
multi_7x28 multi_7x28_mod_8496(clk,rst,matrix_A[8496],matrix_B[96],mul_res1[8496]);
multi_7x28 multi_7x28_mod_8497(clk,rst,matrix_A[8497],matrix_B[97],mul_res1[8497]);
multi_7x28 multi_7x28_mod_8498(clk,rst,matrix_A[8498],matrix_B[98],mul_res1[8498]);
multi_7x28 multi_7x28_mod_8499(clk,rst,matrix_A[8499],matrix_B[99],mul_res1[8499]);
multi_7x28 multi_7x28_mod_8500(clk,rst,matrix_A[8500],matrix_B[100],mul_res1[8500]);
multi_7x28 multi_7x28_mod_8501(clk,rst,matrix_A[8501],matrix_B[101],mul_res1[8501]);
multi_7x28 multi_7x28_mod_8502(clk,rst,matrix_A[8502],matrix_B[102],mul_res1[8502]);
multi_7x28 multi_7x28_mod_8503(clk,rst,matrix_A[8503],matrix_B[103],mul_res1[8503]);
multi_7x28 multi_7x28_mod_8504(clk,rst,matrix_A[8504],matrix_B[104],mul_res1[8504]);
multi_7x28 multi_7x28_mod_8505(clk,rst,matrix_A[8505],matrix_B[105],mul_res1[8505]);
multi_7x28 multi_7x28_mod_8506(clk,rst,matrix_A[8506],matrix_B[106],mul_res1[8506]);
multi_7x28 multi_7x28_mod_8507(clk,rst,matrix_A[8507],matrix_B[107],mul_res1[8507]);
multi_7x28 multi_7x28_mod_8508(clk,rst,matrix_A[8508],matrix_B[108],mul_res1[8508]);
multi_7x28 multi_7x28_mod_8509(clk,rst,matrix_A[8509],matrix_B[109],mul_res1[8509]);
multi_7x28 multi_7x28_mod_8510(clk,rst,matrix_A[8510],matrix_B[110],mul_res1[8510]);
multi_7x28 multi_7x28_mod_8511(clk,rst,matrix_A[8511],matrix_B[111],mul_res1[8511]);
multi_7x28 multi_7x28_mod_8512(clk,rst,matrix_A[8512],matrix_B[112],mul_res1[8512]);
multi_7x28 multi_7x28_mod_8513(clk,rst,matrix_A[8513],matrix_B[113],mul_res1[8513]);
multi_7x28 multi_7x28_mod_8514(clk,rst,matrix_A[8514],matrix_B[114],mul_res1[8514]);
multi_7x28 multi_7x28_mod_8515(clk,rst,matrix_A[8515],matrix_B[115],mul_res1[8515]);
multi_7x28 multi_7x28_mod_8516(clk,rst,matrix_A[8516],matrix_B[116],mul_res1[8516]);
multi_7x28 multi_7x28_mod_8517(clk,rst,matrix_A[8517],matrix_B[117],mul_res1[8517]);
multi_7x28 multi_7x28_mod_8518(clk,rst,matrix_A[8518],matrix_B[118],mul_res1[8518]);
multi_7x28 multi_7x28_mod_8519(clk,rst,matrix_A[8519],matrix_B[119],mul_res1[8519]);
multi_7x28 multi_7x28_mod_8520(clk,rst,matrix_A[8520],matrix_B[120],mul_res1[8520]);
multi_7x28 multi_7x28_mod_8521(clk,rst,matrix_A[8521],matrix_B[121],mul_res1[8521]);
multi_7x28 multi_7x28_mod_8522(clk,rst,matrix_A[8522],matrix_B[122],mul_res1[8522]);
multi_7x28 multi_7x28_mod_8523(clk,rst,matrix_A[8523],matrix_B[123],mul_res1[8523]);
multi_7x28 multi_7x28_mod_8524(clk,rst,matrix_A[8524],matrix_B[124],mul_res1[8524]);
multi_7x28 multi_7x28_mod_8525(clk,rst,matrix_A[8525],matrix_B[125],mul_res1[8525]);
multi_7x28 multi_7x28_mod_8526(clk,rst,matrix_A[8526],matrix_B[126],mul_res1[8526]);
multi_7x28 multi_7x28_mod_8527(clk,rst,matrix_A[8527],matrix_B[127],mul_res1[8527]);
multi_7x28 multi_7x28_mod_8528(clk,rst,matrix_A[8528],matrix_B[128],mul_res1[8528]);
multi_7x28 multi_7x28_mod_8529(clk,rst,matrix_A[8529],matrix_B[129],mul_res1[8529]);
multi_7x28 multi_7x28_mod_8530(clk,rst,matrix_A[8530],matrix_B[130],mul_res1[8530]);
multi_7x28 multi_7x28_mod_8531(clk,rst,matrix_A[8531],matrix_B[131],mul_res1[8531]);
multi_7x28 multi_7x28_mod_8532(clk,rst,matrix_A[8532],matrix_B[132],mul_res1[8532]);
multi_7x28 multi_7x28_mod_8533(clk,rst,matrix_A[8533],matrix_B[133],mul_res1[8533]);
multi_7x28 multi_7x28_mod_8534(clk,rst,matrix_A[8534],matrix_B[134],mul_res1[8534]);
multi_7x28 multi_7x28_mod_8535(clk,rst,matrix_A[8535],matrix_B[135],mul_res1[8535]);
multi_7x28 multi_7x28_mod_8536(clk,rst,matrix_A[8536],matrix_B[136],mul_res1[8536]);
multi_7x28 multi_7x28_mod_8537(clk,rst,matrix_A[8537],matrix_B[137],mul_res1[8537]);
multi_7x28 multi_7x28_mod_8538(clk,rst,matrix_A[8538],matrix_B[138],mul_res1[8538]);
multi_7x28 multi_7x28_mod_8539(clk,rst,matrix_A[8539],matrix_B[139],mul_res1[8539]);
multi_7x28 multi_7x28_mod_8540(clk,rst,matrix_A[8540],matrix_B[140],mul_res1[8540]);
multi_7x28 multi_7x28_mod_8541(clk,rst,matrix_A[8541],matrix_B[141],mul_res1[8541]);
multi_7x28 multi_7x28_mod_8542(clk,rst,matrix_A[8542],matrix_B[142],mul_res1[8542]);
multi_7x28 multi_7x28_mod_8543(clk,rst,matrix_A[8543],matrix_B[143],mul_res1[8543]);
multi_7x28 multi_7x28_mod_8544(clk,rst,matrix_A[8544],matrix_B[144],mul_res1[8544]);
multi_7x28 multi_7x28_mod_8545(clk,rst,matrix_A[8545],matrix_B[145],mul_res1[8545]);
multi_7x28 multi_7x28_mod_8546(clk,rst,matrix_A[8546],matrix_B[146],mul_res1[8546]);
multi_7x28 multi_7x28_mod_8547(clk,rst,matrix_A[8547],matrix_B[147],mul_res1[8547]);
multi_7x28 multi_7x28_mod_8548(clk,rst,matrix_A[8548],matrix_B[148],mul_res1[8548]);
multi_7x28 multi_7x28_mod_8549(clk,rst,matrix_A[8549],matrix_B[149],mul_res1[8549]);
multi_7x28 multi_7x28_mod_8550(clk,rst,matrix_A[8550],matrix_B[150],mul_res1[8550]);
multi_7x28 multi_7x28_mod_8551(clk,rst,matrix_A[8551],matrix_B[151],mul_res1[8551]);
multi_7x28 multi_7x28_mod_8552(clk,rst,matrix_A[8552],matrix_B[152],mul_res1[8552]);
multi_7x28 multi_7x28_mod_8553(clk,rst,matrix_A[8553],matrix_B[153],mul_res1[8553]);
multi_7x28 multi_7x28_mod_8554(clk,rst,matrix_A[8554],matrix_B[154],mul_res1[8554]);
multi_7x28 multi_7x28_mod_8555(clk,rst,matrix_A[8555],matrix_B[155],mul_res1[8555]);
multi_7x28 multi_7x28_mod_8556(clk,rst,matrix_A[8556],matrix_B[156],mul_res1[8556]);
multi_7x28 multi_7x28_mod_8557(clk,rst,matrix_A[8557],matrix_B[157],mul_res1[8557]);
multi_7x28 multi_7x28_mod_8558(clk,rst,matrix_A[8558],matrix_B[158],mul_res1[8558]);
multi_7x28 multi_7x28_mod_8559(clk,rst,matrix_A[8559],matrix_B[159],mul_res1[8559]);
multi_7x28 multi_7x28_mod_8560(clk,rst,matrix_A[8560],matrix_B[160],mul_res1[8560]);
multi_7x28 multi_7x28_mod_8561(clk,rst,matrix_A[8561],matrix_B[161],mul_res1[8561]);
multi_7x28 multi_7x28_mod_8562(clk,rst,matrix_A[8562],matrix_B[162],mul_res1[8562]);
multi_7x28 multi_7x28_mod_8563(clk,rst,matrix_A[8563],matrix_B[163],mul_res1[8563]);
multi_7x28 multi_7x28_mod_8564(clk,rst,matrix_A[8564],matrix_B[164],mul_res1[8564]);
multi_7x28 multi_7x28_mod_8565(clk,rst,matrix_A[8565],matrix_B[165],mul_res1[8565]);
multi_7x28 multi_7x28_mod_8566(clk,rst,matrix_A[8566],matrix_B[166],mul_res1[8566]);
multi_7x28 multi_7x28_mod_8567(clk,rst,matrix_A[8567],matrix_B[167],mul_res1[8567]);
multi_7x28 multi_7x28_mod_8568(clk,rst,matrix_A[8568],matrix_B[168],mul_res1[8568]);
multi_7x28 multi_7x28_mod_8569(clk,rst,matrix_A[8569],matrix_B[169],mul_res1[8569]);
multi_7x28 multi_7x28_mod_8570(clk,rst,matrix_A[8570],matrix_B[170],mul_res1[8570]);
multi_7x28 multi_7x28_mod_8571(clk,rst,matrix_A[8571],matrix_B[171],mul_res1[8571]);
multi_7x28 multi_7x28_mod_8572(clk,rst,matrix_A[8572],matrix_B[172],mul_res1[8572]);
multi_7x28 multi_7x28_mod_8573(clk,rst,matrix_A[8573],matrix_B[173],mul_res1[8573]);
multi_7x28 multi_7x28_mod_8574(clk,rst,matrix_A[8574],matrix_B[174],mul_res1[8574]);
multi_7x28 multi_7x28_mod_8575(clk,rst,matrix_A[8575],matrix_B[175],mul_res1[8575]);
multi_7x28 multi_7x28_mod_8576(clk,rst,matrix_A[8576],matrix_B[176],mul_res1[8576]);
multi_7x28 multi_7x28_mod_8577(clk,rst,matrix_A[8577],matrix_B[177],mul_res1[8577]);
multi_7x28 multi_7x28_mod_8578(clk,rst,matrix_A[8578],matrix_B[178],mul_res1[8578]);
multi_7x28 multi_7x28_mod_8579(clk,rst,matrix_A[8579],matrix_B[179],mul_res1[8579]);
multi_7x28 multi_7x28_mod_8580(clk,rst,matrix_A[8580],matrix_B[180],mul_res1[8580]);
multi_7x28 multi_7x28_mod_8581(clk,rst,matrix_A[8581],matrix_B[181],mul_res1[8581]);
multi_7x28 multi_7x28_mod_8582(clk,rst,matrix_A[8582],matrix_B[182],mul_res1[8582]);
multi_7x28 multi_7x28_mod_8583(clk,rst,matrix_A[8583],matrix_B[183],mul_res1[8583]);
multi_7x28 multi_7x28_mod_8584(clk,rst,matrix_A[8584],matrix_B[184],mul_res1[8584]);
multi_7x28 multi_7x28_mod_8585(clk,rst,matrix_A[8585],matrix_B[185],mul_res1[8585]);
multi_7x28 multi_7x28_mod_8586(clk,rst,matrix_A[8586],matrix_B[186],mul_res1[8586]);
multi_7x28 multi_7x28_mod_8587(clk,rst,matrix_A[8587],matrix_B[187],mul_res1[8587]);
multi_7x28 multi_7x28_mod_8588(clk,rst,matrix_A[8588],matrix_B[188],mul_res1[8588]);
multi_7x28 multi_7x28_mod_8589(clk,rst,matrix_A[8589],matrix_B[189],mul_res1[8589]);
multi_7x28 multi_7x28_mod_8590(clk,rst,matrix_A[8590],matrix_B[190],mul_res1[8590]);
multi_7x28 multi_7x28_mod_8591(clk,rst,matrix_A[8591],matrix_B[191],mul_res1[8591]);
multi_7x28 multi_7x28_mod_8592(clk,rst,matrix_A[8592],matrix_B[192],mul_res1[8592]);
multi_7x28 multi_7x28_mod_8593(clk,rst,matrix_A[8593],matrix_B[193],mul_res1[8593]);
multi_7x28 multi_7x28_mod_8594(clk,rst,matrix_A[8594],matrix_B[194],mul_res1[8594]);
multi_7x28 multi_7x28_mod_8595(clk,rst,matrix_A[8595],matrix_B[195],mul_res1[8595]);
multi_7x28 multi_7x28_mod_8596(clk,rst,matrix_A[8596],matrix_B[196],mul_res1[8596]);
multi_7x28 multi_7x28_mod_8597(clk,rst,matrix_A[8597],matrix_B[197],mul_res1[8597]);
multi_7x28 multi_7x28_mod_8598(clk,rst,matrix_A[8598],matrix_B[198],mul_res1[8598]);
multi_7x28 multi_7x28_mod_8599(clk,rst,matrix_A[8599],matrix_B[199],mul_res1[8599]);
multi_7x28 multi_7x28_mod_8600(clk,rst,matrix_A[8600],matrix_B[0],mul_res1[8600]);
multi_7x28 multi_7x28_mod_8601(clk,rst,matrix_A[8601],matrix_B[1],mul_res1[8601]);
multi_7x28 multi_7x28_mod_8602(clk,rst,matrix_A[8602],matrix_B[2],mul_res1[8602]);
multi_7x28 multi_7x28_mod_8603(clk,rst,matrix_A[8603],matrix_B[3],mul_res1[8603]);
multi_7x28 multi_7x28_mod_8604(clk,rst,matrix_A[8604],matrix_B[4],mul_res1[8604]);
multi_7x28 multi_7x28_mod_8605(clk,rst,matrix_A[8605],matrix_B[5],mul_res1[8605]);
multi_7x28 multi_7x28_mod_8606(clk,rst,matrix_A[8606],matrix_B[6],mul_res1[8606]);
multi_7x28 multi_7x28_mod_8607(clk,rst,matrix_A[8607],matrix_B[7],mul_res1[8607]);
multi_7x28 multi_7x28_mod_8608(clk,rst,matrix_A[8608],matrix_B[8],mul_res1[8608]);
multi_7x28 multi_7x28_mod_8609(clk,rst,matrix_A[8609],matrix_B[9],mul_res1[8609]);
multi_7x28 multi_7x28_mod_8610(clk,rst,matrix_A[8610],matrix_B[10],mul_res1[8610]);
multi_7x28 multi_7x28_mod_8611(clk,rst,matrix_A[8611],matrix_B[11],mul_res1[8611]);
multi_7x28 multi_7x28_mod_8612(clk,rst,matrix_A[8612],matrix_B[12],mul_res1[8612]);
multi_7x28 multi_7x28_mod_8613(clk,rst,matrix_A[8613],matrix_B[13],mul_res1[8613]);
multi_7x28 multi_7x28_mod_8614(clk,rst,matrix_A[8614],matrix_B[14],mul_res1[8614]);
multi_7x28 multi_7x28_mod_8615(clk,rst,matrix_A[8615],matrix_B[15],mul_res1[8615]);
multi_7x28 multi_7x28_mod_8616(clk,rst,matrix_A[8616],matrix_B[16],mul_res1[8616]);
multi_7x28 multi_7x28_mod_8617(clk,rst,matrix_A[8617],matrix_B[17],mul_res1[8617]);
multi_7x28 multi_7x28_mod_8618(clk,rst,matrix_A[8618],matrix_B[18],mul_res1[8618]);
multi_7x28 multi_7x28_mod_8619(clk,rst,matrix_A[8619],matrix_B[19],mul_res1[8619]);
multi_7x28 multi_7x28_mod_8620(clk,rst,matrix_A[8620],matrix_B[20],mul_res1[8620]);
multi_7x28 multi_7x28_mod_8621(clk,rst,matrix_A[8621],matrix_B[21],mul_res1[8621]);
multi_7x28 multi_7x28_mod_8622(clk,rst,matrix_A[8622],matrix_B[22],mul_res1[8622]);
multi_7x28 multi_7x28_mod_8623(clk,rst,matrix_A[8623],matrix_B[23],mul_res1[8623]);
multi_7x28 multi_7x28_mod_8624(clk,rst,matrix_A[8624],matrix_B[24],mul_res1[8624]);
multi_7x28 multi_7x28_mod_8625(clk,rst,matrix_A[8625],matrix_B[25],mul_res1[8625]);
multi_7x28 multi_7x28_mod_8626(clk,rst,matrix_A[8626],matrix_B[26],mul_res1[8626]);
multi_7x28 multi_7x28_mod_8627(clk,rst,matrix_A[8627],matrix_B[27],mul_res1[8627]);
multi_7x28 multi_7x28_mod_8628(clk,rst,matrix_A[8628],matrix_B[28],mul_res1[8628]);
multi_7x28 multi_7x28_mod_8629(clk,rst,matrix_A[8629],matrix_B[29],mul_res1[8629]);
multi_7x28 multi_7x28_mod_8630(clk,rst,matrix_A[8630],matrix_B[30],mul_res1[8630]);
multi_7x28 multi_7x28_mod_8631(clk,rst,matrix_A[8631],matrix_B[31],mul_res1[8631]);
multi_7x28 multi_7x28_mod_8632(clk,rst,matrix_A[8632],matrix_B[32],mul_res1[8632]);
multi_7x28 multi_7x28_mod_8633(clk,rst,matrix_A[8633],matrix_B[33],mul_res1[8633]);
multi_7x28 multi_7x28_mod_8634(clk,rst,matrix_A[8634],matrix_B[34],mul_res1[8634]);
multi_7x28 multi_7x28_mod_8635(clk,rst,matrix_A[8635],matrix_B[35],mul_res1[8635]);
multi_7x28 multi_7x28_mod_8636(clk,rst,matrix_A[8636],matrix_B[36],mul_res1[8636]);
multi_7x28 multi_7x28_mod_8637(clk,rst,matrix_A[8637],matrix_B[37],mul_res1[8637]);
multi_7x28 multi_7x28_mod_8638(clk,rst,matrix_A[8638],matrix_B[38],mul_res1[8638]);
multi_7x28 multi_7x28_mod_8639(clk,rst,matrix_A[8639],matrix_B[39],mul_res1[8639]);
multi_7x28 multi_7x28_mod_8640(clk,rst,matrix_A[8640],matrix_B[40],mul_res1[8640]);
multi_7x28 multi_7x28_mod_8641(clk,rst,matrix_A[8641],matrix_B[41],mul_res1[8641]);
multi_7x28 multi_7x28_mod_8642(clk,rst,matrix_A[8642],matrix_B[42],mul_res1[8642]);
multi_7x28 multi_7x28_mod_8643(clk,rst,matrix_A[8643],matrix_B[43],mul_res1[8643]);
multi_7x28 multi_7x28_mod_8644(clk,rst,matrix_A[8644],matrix_B[44],mul_res1[8644]);
multi_7x28 multi_7x28_mod_8645(clk,rst,matrix_A[8645],matrix_B[45],mul_res1[8645]);
multi_7x28 multi_7x28_mod_8646(clk,rst,matrix_A[8646],matrix_B[46],mul_res1[8646]);
multi_7x28 multi_7x28_mod_8647(clk,rst,matrix_A[8647],matrix_B[47],mul_res1[8647]);
multi_7x28 multi_7x28_mod_8648(clk,rst,matrix_A[8648],matrix_B[48],mul_res1[8648]);
multi_7x28 multi_7x28_mod_8649(clk,rst,matrix_A[8649],matrix_B[49],mul_res1[8649]);
multi_7x28 multi_7x28_mod_8650(clk,rst,matrix_A[8650],matrix_B[50],mul_res1[8650]);
multi_7x28 multi_7x28_mod_8651(clk,rst,matrix_A[8651],matrix_B[51],mul_res1[8651]);
multi_7x28 multi_7x28_mod_8652(clk,rst,matrix_A[8652],matrix_B[52],mul_res1[8652]);
multi_7x28 multi_7x28_mod_8653(clk,rst,matrix_A[8653],matrix_B[53],mul_res1[8653]);
multi_7x28 multi_7x28_mod_8654(clk,rst,matrix_A[8654],matrix_B[54],mul_res1[8654]);
multi_7x28 multi_7x28_mod_8655(clk,rst,matrix_A[8655],matrix_B[55],mul_res1[8655]);
multi_7x28 multi_7x28_mod_8656(clk,rst,matrix_A[8656],matrix_B[56],mul_res1[8656]);
multi_7x28 multi_7x28_mod_8657(clk,rst,matrix_A[8657],matrix_B[57],mul_res1[8657]);
multi_7x28 multi_7x28_mod_8658(clk,rst,matrix_A[8658],matrix_B[58],mul_res1[8658]);
multi_7x28 multi_7x28_mod_8659(clk,rst,matrix_A[8659],matrix_B[59],mul_res1[8659]);
multi_7x28 multi_7x28_mod_8660(clk,rst,matrix_A[8660],matrix_B[60],mul_res1[8660]);
multi_7x28 multi_7x28_mod_8661(clk,rst,matrix_A[8661],matrix_B[61],mul_res1[8661]);
multi_7x28 multi_7x28_mod_8662(clk,rst,matrix_A[8662],matrix_B[62],mul_res1[8662]);
multi_7x28 multi_7x28_mod_8663(clk,rst,matrix_A[8663],matrix_B[63],mul_res1[8663]);
multi_7x28 multi_7x28_mod_8664(clk,rst,matrix_A[8664],matrix_B[64],mul_res1[8664]);
multi_7x28 multi_7x28_mod_8665(clk,rst,matrix_A[8665],matrix_B[65],mul_res1[8665]);
multi_7x28 multi_7x28_mod_8666(clk,rst,matrix_A[8666],matrix_B[66],mul_res1[8666]);
multi_7x28 multi_7x28_mod_8667(clk,rst,matrix_A[8667],matrix_B[67],mul_res1[8667]);
multi_7x28 multi_7x28_mod_8668(clk,rst,matrix_A[8668],matrix_B[68],mul_res1[8668]);
multi_7x28 multi_7x28_mod_8669(clk,rst,matrix_A[8669],matrix_B[69],mul_res1[8669]);
multi_7x28 multi_7x28_mod_8670(clk,rst,matrix_A[8670],matrix_B[70],mul_res1[8670]);
multi_7x28 multi_7x28_mod_8671(clk,rst,matrix_A[8671],matrix_B[71],mul_res1[8671]);
multi_7x28 multi_7x28_mod_8672(clk,rst,matrix_A[8672],matrix_B[72],mul_res1[8672]);
multi_7x28 multi_7x28_mod_8673(clk,rst,matrix_A[8673],matrix_B[73],mul_res1[8673]);
multi_7x28 multi_7x28_mod_8674(clk,rst,matrix_A[8674],matrix_B[74],mul_res1[8674]);
multi_7x28 multi_7x28_mod_8675(clk,rst,matrix_A[8675],matrix_B[75],mul_res1[8675]);
multi_7x28 multi_7x28_mod_8676(clk,rst,matrix_A[8676],matrix_B[76],mul_res1[8676]);
multi_7x28 multi_7x28_mod_8677(clk,rst,matrix_A[8677],matrix_B[77],mul_res1[8677]);
multi_7x28 multi_7x28_mod_8678(clk,rst,matrix_A[8678],matrix_B[78],mul_res1[8678]);
multi_7x28 multi_7x28_mod_8679(clk,rst,matrix_A[8679],matrix_B[79],mul_res1[8679]);
multi_7x28 multi_7x28_mod_8680(clk,rst,matrix_A[8680],matrix_B[80],mul_res1[8680]);
multi_7x28 multi_7x28_mod_8681(clk,rst,matrix_A[8681],matrix_B[81],mul_res1[8681]);
multi_7x28 multi_7x28_mod_8682(clk,rst,matrix_A[8682],matrix_B[82],mul_res1[8682]);
multi_7x28 multi_7x28_mod_8683(clk,rst,matrix_A[8683],matrix_B[83],mul_res1[8683]);
multi_7x28 multi_7x28_mod_8684(clk,rst,matrix_A[8684],matrix_B[84],mul_res1[8684]);
multi_7x28 multi_7x28_mod_8685(clk,rst,matrix_A[8685],matrix_B[85],mul_res1[8685]);
multi_7x28 multi_7x28_mod_8686(clk,rst,matrix_A[8686],matrix_B[86],mul_res1[8686]);
multi_7x28 multi_7x28_mod_8687(clk,rst,matrix_A[8687],matrix_B[87],mul_res1[8687]);
multi_7x28 multi_7x28_mod_8688(clk,rst,matrix_A[8688],matrix_B[88],mul_res1[8688]);
multi_7x28 multi_7x28_mod_8689(clk,rst,matrix_A[8689],matrix_B[89],mul_res1[8689]);
multi_7x28 multi_7x28_mod_8690(clk,rst,matrix_A[8690],matrix_B[90],mul_res1[8690]);
multi_7x28 multi_7x28_mod_8691(clk,rst,matrix_A[8691],matrix_B[91],mul_res1[8691]);
multi_7x28 multi_7x28_mod_8692(clk,rst,matrix_A[8692],matrix_B[92],mul_res1[8692]);
multi_7x28 multi_7x28_mod_8693(clk,rst,matrix_A[8693],matrix_B[93],mul_res1[8693]);
multi_7x28 multi_7x28_mod_8694(clk,rst,matrix_A[8694],matrix_B[94],mul_res1[8694]);
multi_7x28 multi_7x28_mod_8695(clk,rst,matrix_A[8695],matrix_B[95],mul_res1[8695]);
multi_7x28 multi_7x28_mod_8696(clk,rst,matrix_A[8696],matrix_B[96],mul_res1[8696]);
multi_7x28 multi_7x28_mod_8697(clk,rst,matrix_A[8697],matrix_B[97],mul_res1[8697]);
multi_7x28 multi_7x28_mod_8698(clk,rst,matrix_A[8698],matrix_B[98],mul_res1[8698]);
multi_7x28 multi_7x28_mod_8699(clk,rst,matrix_A[8699],matrix_B[99],mul_res1[8699]);
multi_7x28 multi_7x28_mod_8700(clk,rst,matrix_A[8700],matrix_B[100],mul_res1[8700]);
multi_7x28 multi_7x28_mod_8701(clk,rst,matrix_A[8701],matrix_B[101],mul_res1[8701]);
multi_7x28 multi_7x28_mod_8702(clk,rst,matrix_A[8702],matrix_B[102],mul_res1[8702]);
multi_7x28 multi_7x28_mod_8703(clk,rst,matrix_A[8703],matrix_B[103],mul_res1[8703]);
multi_7x28 multi_7x28_mod_8704(clk,rst,matrix_A[8704],matrix_B[104],mul_res1[8704]);
multi_7x28 multi_7x28_mod_8705(clk,rst,matrix_A[8705],matrix_B[105],mul_res1[8705]);
multi_7x28 multi_7x28_mod_8706(clk,rst,matrix_A[8706],matrix_B[106],mul_res1[8706]);
multi_7x28 multi_7x28_mod_8707(clk,rst,matrix_A[8707],matrix_B[107],mul_res1[8707]);
multi_7x28 multi_7x28_mod_8708(clk,rst,matrix_A[8708],matrix_B[108],mul_res1[8708]);
multi_7x28 multi_7x28_mod_8709(clk,rst,matrix_A[8709],matrix_B[109],mul_res1[8709]);
multi_7x28 multi_7x28_mod_8710(clk,rst,matrix_A[8710],matrix_B[110],mul_res1[8710]);
multi_7x28 multi_7x28_mod_8711(clk,rst,matrix_A[8711],matrix_B[111],mul_res1[8711]);
multi_7x28 multi_7x28_mod_8712(clk,rst,matrix_A[8712],matrix_B[112],mul_res1[8712]);
multi_7x28 multi_7x28_mod_8713(clk,rst,matrix_A[8713],matrix_B[113],mul_res1[8713]);
multi_7x28 multi_7x28_mod_8714(clk,rst,matrix_A[8714],matrix_B[114],mul_res1[8714]);
multi_7x28 multi_7x28_mod_8715(clk,rst,matrix_A[8715],matrix_B[115],mul_res1[8715]);
multi_7x28 multi_7x28_mod_8716(clk,rst,matrix_A[8716],matrix_B[116],mul_res1[8716]);
multi_7x28 multi_7x28_mod_8717(clk,rst,matrix_A[8717],matrix_B[117],mul_res1[8717]);
multi_7x28 multi_7x28_mod_8718(clk,rst,matrix_A[8718],matrix_B[118],mul_res1[8718]);
multi_7x28 multi_7x28_mod_8719(clk,rst,matrix_A[8719],matrix_B[119],mul_res1[8719]);
multi_7x28 multi_7x28_mod_8720(clk,rst,matrix_A[8720],matrix_B[120],mul_res1[8720]);
multi_7x28 multi_7x28_mod_8721(clk,rst,matrix_A[8721],matrix_B[121],mul_res1[8721]);
multi_7x28 multi_7x28_mod_8722(clk,rst,matrix_A[8722],matrix_B[122],mul_res1[8722]);
multi_7x28 multi_7x28_mod_8723(clk,rst,matrix_A[8723],matrix_B[123],mul_res1[8723]);
multi_7x28 multi_7x28_mod_8724(clk,rst,matrix_A[8724],matrix_B[124],mul_res1[8724]);
multi_7x28 multi_7x28_mod_8725(clk,rst,matrix_A[8725],matrix_B[125],mul_res1[8725]);
multi_7x28 multi_7x28_mod_8726(clk,rst,matrix_A[8726],matrix_B[126],mul_res1[8726]);
multi_7x28 multi_7x28_mod_8727(clk,rst,matrix_A[8727],matrix_B[127],mul_res1[8727]);
multi_7x28 multi_7x28_mod_8728(clk,rst,matrix_A[8728],matrix_B[128],mul_res1[8728]);
multi_7x28 multi_7x28_mod_8729(clk,rst,matrix_A[8729],matrix_B[129],mul_res1[8729]);
multi_7x28 multi_7x28_mod_8730(clk,rst,matrix_A[8730],matrix_B[130],mul_res1[8730]);
multi_7x28 multi_7x28_mod_8731(clk,rst,matrix_A[8731],matrix_B[131],mul_res1[8731]);
multi_7x28 multi_7x28_mod_8732(clk,rst,matrix_A[8732],matrix_B[132],mul_res1[8732]);
multi_7x28 multi_7x28_mod_8733(clk,rst,matrix_A[8733],matrix_B[133],mul_res1[8733]);
multi_7x28 multi_7x28_mod_8734(clk,rst,matrix_A[8734],matrix_B[134],mul_res1[8734]);
multi_7x28 multi_7x28_mod_8735(clk,rst,matrix_A[8735],matrix_B[135],mul_res1[8735]);
multi_7x28 multi_7x28_mod_8736(clk,rst,matrix_A[8736],matrix_B[136],mul_res1[8736]);
multi_7x28 multi_7x28_mod_8737(clk,rst,matrix_A[8737],matrix_B[137],mul_res1[8737]);
multi_7x28 multi_7x28_mod_8738(clk,rst,matrix_A[8738],matrix_B[138],mul_res1[8738]);
multi_7x28 multi_7x28_mod_8739(clk,rst,matrix_A[8739],matrix_B[139],mul_res1[8739]);
multi_7x28 multi_7x28_mod_8740(clk,rst,matrix_A[8740],matrix_B[140],mul_res1[8740]);
multi_7x28 multi_7x28_mod_8741(clk,rst,matrix_A[8741],matrix_B[141],mul_res1[8741]);
multi_7x28 multi_7x28_mod_8742(clk,rst,matrix_A[8742],matrix_B[142],mul_res1[8742]);
multi_7x28 multi_7x28_mod_8743(clk,rst,matrix_A[8743],matrix_B[143],mul_res1[8743]);
multi_7x28 multi_7x28_mod_8744(clk,rst,matrix_A[8744],matrix_B[144],mul_res1[8744]);
multi_7x28 multi_7x28_mod_8745(clk,rst,matrix_A[8745],matrix_B[145],mul_res1[8745]);
multi_7x28 multi_7x28_mod_8746(clk,rst,matrix_A[8746],matrix_B[146],mul_res1[8746]);
multi_7x28 multi_7x28_mod_8747(clk,rst,matrix_A[8747],matrix_B[147],mul_res1[8747]);
multi_7x28 multi_7x28_mod_8748(clk,rst,matrix_A[8748],matrix_B[148],mul_res1[8748]);
multi_7x28 multi_7x28_mod_8749(clk,rst,matrix_A[8749],matrix_B[149],mul_res1[8749]);
multi_7x28 multi_7x28_mod_8750(clk,rst,matrix_A[8750],matrix_B[150],mul_res1[8750]);
multi_7x28 multi_7x28_mod_8751(clk,rst,matrix_A[8751],matrix_B[151],mul_res1[8751]);
multi_7x28 multi_7x28_mod_8752(clk,rst,matrix_A[8752],matrix_B[152],mul_res1[8752]);
multi_7x28 multi_7x28_mod_8753(clk,rst,matrix_A[8753],matrix_B[153],mul_res1[8753]);
multi_7x28 multi_7x28_mod_8754(clk,rst,matrix_A[8754],matrix_B[154],mul_res1[8754]);
multi_7x28 multi_7x28_mod_8755(clk,rst,matrix_A[8755],matrix_B[155],mul_res1[8755]);
multi_7x28 multi_7x28_mod_8756(clk,rst,matrix_A[8756],matrix_B[156],mul_res1[8756]);
multi_7x28 multi_7x28_mod_8757(clk,rst,matrix_A[8757],matrix_B[157],mul_res1[8757]);
multi_7x28 multi_7x28_mod_8758(clk,rst,matrix_A[8758],matrix_B[158],mul_res1[8758]);
multi_7x28 multi_7x28_mod_8759(clk,rst,matrix_A[8759],matrix_B[159],mul_res1[8759]);
multi_7x28 multi_7x28_mod_8760(clk,rst,matrix_A[8760],matrix_B[160],mul_res1[8760]);
multi_7x28 multi_7x28_mod_8761(clk,rst,matrix_A[8761],matrix_B[161],mul_res1[8761]);
multi_7x28 multi_7x28_mod_8762(clk,rst,matrix_A[8762],matrix_B[162],mul_res1[8762]);
multi_7x28 multi_7x28_mod_8763(clk,rst,matrix_A[8763],matrix_B[163],mul_res1[8763]);
multi_7x28 multi_7x28_mod_8764(clk,rst,matrix_A[8764],matrix_B[164],mul_res1[8764]);
multi_7x28 multi_7x28_mod_8765(clk,rst,matrix_A[8765],matrix_B[165],mul_res1[8765]);
multi_7x28 multi_7x28_mod_8766(clk,rst,matrix_A[8766],matrix_B[166],mul_res1[8766]);
multi_7x28 multi_7x28_mod_8767(clk,rst,matrix_A[8767],matrix_B[167],mul_res1[8767]);
multi_7x28 multi_7x28_mod_8768(clk,rst,matrix_A[8768],matrix_B[168],mul_res1[8768]);
multi_7x28 multi_7x28_mod_8769(clk,rst,matrix_A[8769],matrix_B[169],mul_res1[8769]);
multi_7x28 multi_7x28_mod_8770(clk,rst,matrix_A[8770],matrix_B[170],mul_res1[8770]);
multi_7x28 multi_7x28_mod_8771(clk,rst,matrix_A[8771],matrix_B[171],mul_res1[8771]);
multi_7x28 multi_7x28_mod_8772(clk,rst,matrix_A[8772],matrix_B[172],mul_res1[8772]);
multi_7x28 multi_7x28_mod_8773(clk,rst,matrix_A[8773],matrix_B[173],mul_res1[8773]);
multi_7x28 multi_7x28_mod_8774(clk,rst,matrix_A[8774],matrix_B[174],mul_res1[8774]);
multi_7x28 multi_7x28_mod_8775(clk,rst,matrix_A[8775],matrix_B[175],mul_res1[8775]);
multi_7x28 multi_7x28_mod_8776(clk,rst,matrix_A[8776],matrix_B[176],mul_res1[8776]);
multi_7x28 multi_7x28_mod_8777(clk,rst,matrix_A[8777],matrix_B[177],mul_res1[8777]);
multi_7x28 multi_7x28_mod_8778(clk,rst,matrix_A[8778],matrix_B[178],mul_res1[8778]);
multi_7x28 multi_7x28_mod_8779(clk,rst,matrix_A[8779],matrix_B[179],mul_res1[8779]);
multi_7x28 multi_7x28_mod_8780(clk,rst,matrix_A[8780],matrix_B[180],mul_res1[8780]);
multi_7x28 multi_7x28_mod_8781(clk,rst,matrix_A[8781],matrix_B[181],mul_res1[8781]);
multi_7x28 multi_7x28_mod_8782(clk,rst,matrix_A[8782],matrix_B[182],mul_res1[8782]);
multi_7x28 multi_7x28_mod_8783(clk,rst,matrix_A[8783],matrix_B[183],mul_res1[8783]);
multi_7x28 multi_7x28_mod_8784(clk,rst,matrix_A[8784],matrix_B[184],mul_res1[8784]);
multi_7x28 multi_7x28_mod_8785(clk,rst,matrix_A[8785],matrix_B[185],mul_res1[8785]);
multi_7x28 multi_7x28_mod_8786(clk,rst,matrix_A[8786],matrix_B[186],mul_res1[8786]);
multi_7x28 multi_7x28_mod_8787(clk,rst,matrix_A[8787],matrix_B[187],mul_res1[8787]);
multi_7x28 multi_7x28_mod_8788(clk,rst,matrix_A[8788],matrix_B[188],mul_res1[8788]);
multi_7x28 multi_7x28_mod_8789(clk,rst,matrix_A[8789],matrix_B[189],mul_res1[8789]);
multi_7x28 multi_7x28_mod_8790(clk,rst,matrix_A[8790],matrix_B[190],mul_res1[8790]);
multi_7x28 multi_7x28_mod_8791(clk,rst,matrix_A[8791],matrix_B[191],mul_res1[8791]);
multi_7x28 multi_7x28_mod_8792(clk,rst,matrix_A[8792],matrix_B[192],mul_res1[8792]);
multi_7x28 multi_7x28_mod_8793(clk,rst,matrix_A[8793],matrix_B[193],mul_res1[8793]);
multi_7x28 multi_7x28_mod_8794(clk,rst,matrix_A[8794],matrix_B[194],mul_res1[8794]);
multi_7x28 multi_7x28_mod_8795(clk,rst,matrix_A[8795],matrix_B[195],mul_res1[8795]);
multi_7x28 multi_7x28_mod_8796(clk,rst,matrix_A[8796],matrix_B[196],mul_res1[8796]);
multi_7x28 multi_7x28_mod_8797(clk,rst,matrix_A[8797],matrix_B[197],mul_res1[8797]);
multi_7x28 multi_7x28_mod_8798(clk,rst,matrix_A[8798],matrix_B[198],mul_res1[8798]);
multi_7x28 multi_7x28_mod_8799(clk,rst,matrix_A[8799],matrix_B[199],mul_res1[8799]);
multi_7x28 multi_7x28_mod_8800(clk,rst,matrix_A[8800],matrix_B[0],mul_res1[8800]);
multi_7x28 multi_7x28_mod_8801(clk,rst,matrix_A[8801],matrix_B[1],mul_res1[8801]);
multi_7x28 multi_7x28_mod_8802(clk,rst,matrix_A[8802],matrix_B[2],mul_res1[8802]);
multi_7x28 multi_7x28_mod_8803(clk,rst,matrix_A[8803],matrix_B[3],mul_res1[8803]);
multi_7x28 multi_7x28_mod_8804(clk,rst,matrix_A[8804],matrix_B[4],mul_res1[8804]);
multi_7x28 multi_7x28_mod_8805(clk,rst,matrix_A[8805],matrix_B[5],mul_res1[8805]);
multi_7x28 multi_7x28_mod_8806(clk,rst,matrix_A[8806],matrix_B[6],mul_res1[8806]);
multi_7x28 multi_7x28_mod_8807(clk,rst,matrix_A[8807],matrix_B[7],mul_res1[8807]);
multi_7x28 multi_7x28_mod_8808(clk,rst,matrix_A[8808],matrix_B[8],mul_res1[8808]);
multi_7x28 multi_7x28_mod_8809(clk,rst,matrix_A[8809],matrix_B[9],mul_res1[8809]);
multi_7x28 multi_7x28_mod_8810(clk,rst,matrix_A[8810],matrix_B[10],mul_res1[8810]);
multi_7x28 multi_7x28_mod_8811(clk,rst,matrix_A[8811],matrix_B[11],mul_res1[8811]);
multi_7x28 multi_7x28_mod_8812(clk,rst,matrix_A[8812],matrix_B[12],mul_res1[8812]);
multi_7x28 multi_7x28_mod_8813(clk,rst,matrix_A[8813],matrix_B[13],mul_res1[8813]);
multi_7x28 multi_7x28_mod_8814(clk,rst,matrix_A[8814],matrix_B[14],mul_res1[8814]);
multi_7x28 multi_7x28_mod_8815(clk,rst,matrix_A[8815],matrix_B[15],mul_res1[8815]);
multi_7x28 multi_7x28_mod_8816(clk,rst,matrix_A[8816],matrix_B[16],mul_res1[8816]);
multi_7x28 multi_7x28_mod_8817(clk,rst,matrix_A[8817],matrix_B[17],mul_res1[8817]);
multi_7x28 multi_7x28_mod_8818(clk,rst,matrix_A[8818],matrix_B[18],mul_res1[8818]);
multi_7x28 multi_7x28_mod_8819(clk,rst,matrix_A[8819],matrix_B[19],mul_res1[8819]);
multi_7x28 multi_7x28_mod_8820(clk,rst,matrix_A[8820],matrix_B[20],mul_res1[8820]);
multi_7x28 multi_7x28_mod_8821(clk,rst,matrix_A[8821],matrix_B[21],mul_res1[8821]);
multi_7x28 multi_7x28_mod_8822(clk,rst,matrix_A[8822],matrix_B[22],mul_res1[8822]);
multi_7x28 multi_7x28_mod_8823(clk,rst,matrix_A[8823],matrix_B[23],mul_res1[8823]);
multi_7x28 multi_7x28_mod_8824(clk,rst,matrix_A[8824],matrix_B[24],mul_res1[8824]);
multi_7x28 multi_7x28_mod_8825(clk,rst,matrix_A[8825],matrix_B[25],mul_res1[8825]);
multi_7x28 multi_7x28_mod_8826(clk,rst,matrix_A[8826],matrix_B[26],mul_res1[8826]);
multi_7x28 multi_7x28_mod_8827(clk,rst,matrix_A[8827],matrix_B[27],mul_res1[8827]);
multi_7x28 multi_7x28_mod_8828(clk,rst,matrix_A[8828],matrix_B[28],mul_res1[8828]);
multi_7x28 multi_7x28_mod_8829(clk,rst,matrix_A[8829],matrix_B[29],mul_res1[8829]);
multi_7x28 multi_7x28_mod_8830(clk,rst,matrix_A[8830],matrix_B[30],mul_res1[8830]);
multi_7x28 multi_7x28_mod_8831(clk,rst,matrix_A[8831],matrix_B[31],mul_res1[8831]);
multi_7x28 multi_7x28_mod_8832(clk,rst,matrix_A[8832],matrix_B[32],mul_res1[8832]);
multi_7x28 multi_7x28_mod_8833(clk,rst,matrix_A[8833],matrix_B[33],mul_res1[8833]);
multi_7x28 multi_7x28_mod_8834(clk,rst,matrix_A[8834],matrix_B[34],mul_res1[8834]);
multi_7x28 multi_7x28_mod_8835(clk,rst,matrix_A[8835],matrix_B[35],mul_res1[8835]);
multi_7x28 multi_7x28_mod_8836(clk,rst,matrix_A[8836],matrix_B[36],mul_res1[8836]);
multi_7x28 multi_7x28_mod_8837(clk,rst,matrix_A[8837],matrix_B[37],mul_res1[8837]);
multi_7x28 multi_7x28_mod_8838(clk,rst,matrix_A[8838],matrix_B[38],mul_res1[8838]);
multi_7x28 multi_7x28_mod_8839(clk,rst,matrix_A[8839],matrix_B[39],mul_res1[8839]);
multi_7x28 multi_7x28_mod_8840(clk,rst,matrix_A[8840],matrix_B[40],mul_res1[8840]);
multi_7x28 multi_7x28_mod_8841(clk,rst,matrix_A[8841],matrix_B[41],mul_res1[8841]);
multi_7x28 multi_7x28_mod_8842(clk,rst,matrix_A[8842],matrix_B[42],mul_res1[8842]);
multi_7x28 multi_7x28_mod_8843(clk,rst,matrix_A[8843],matrix_B[43],mul_res1[8843]);
multi_7x28 multi_7x28_mod_8844(clk,rst,matrix_A[8844],matrix_B[44],mul_res1[8844]);
multi_7x28 multi_7x28_mod_8845(clk,rst,matrix_A[8845],matrix_B[45],mul_res1[8845]);
multi_7x28 multi_7x28_mod_8846(clk,rst,matrix_A[8846],matrix_B[46],mul_res1[8846]);
multi_7x28 multi_7x28_mod_8847(clk,rst,matrix_A[8847],matrix_B[47],mul_res1[8847]);
multi_7x28 multi_7x28_mod_8848(clk,rst,matrix_A[8848],matrix_B[48],mul_res1[8848]);
multi_7x28 multi_7x28_mod_8849(clk,rst,matrix_A[8849],matrix_B[49],mul_res1[8849]);
multi_7x28 multi_7x28_mod_8850(clk,rst,matrix_A[8850],matrix_B[50],mul_res1[8850]);
multi_7x28 multi_7x28_mod_8851(clk,rst,matrix_A[8851],matrix_B[51],mul_res1[8851]);
multi_7x28 multi_7x28_mod_8852(clk,rst,matrix_A[8852],matrix_B[52],mul_res1[8852]);
multi_7x28 multi_7x28_mod_8853(clk,rst,matrix_A[8853],matrix_B[53],mul_res1[8853]);
multi_7x28 multi_7x28_mod_8854(clk,rst,matrix_A[8854],matrix_B[54],mul_res1[8854]);
multi_7x28 multi_7x28_mod_8855(clk,rst,matrix_A[8855],matrix_B[55],mul_res1[8855]);
multi_7x28 multi_7x28_mod_8856(clk,rst,matrix_A[8856],matrix_B[56],mul_res1[8856]);
multi_7x28 multi_7x28_mod_8857(clk,rst,matrix_A[8857],matrix_B[57],mul_res1[8857]);
multi_7x28 multi_7x28_mod_8858(clk,rst,matrix_A[8858],matrix_B[58],mul_res1[8858]);
multi_7x28 multi_7x28_mod_8859(clk,rst,matrix_A[8859],matrix_B[59],mul_res1[8859]);
multi_7x28 multi_7x28_mod_8860(clk,rst,matrix_A[8860],matrix_B[60],mul_res1[8860]);
multi_7x28 multi_7x28_mod_8861(clk,rst,matrix_A[8861],matrix_B[61],mul_res1[8861]);
multi_7x28 multi_7x28_mod_8862(clk,rst,matrix_A[8862],matrix_B[62],mul_res1[8862]);
multi_7x28 multi_7x28_mod_8863(clk,rst,matrix_A[8863],matrix_B[63],mul_res1[8863]);
multi_7x28 multi_7x28_mod_8864(clk,rst,matrix_A[8864],matrix_B[64],mul_res1[8864]);
multi_7x28 multi_7x28_mod_8865(clk,rst,matrix_A[8865],matrix_B[65],mul_res1[8865]);
multi_7x28 multi_7x28_mod_8866(clk,rst,matrix_A[8866],matrix_B[66],mul_res1[8866]);
multi_7x28 multi_7x28_mod_8867(clk,rst,matrix_A[8867],matrix_B[67],mul_res1[8867]);
multi_7x28 multi_7x28_mod_8868(clk,rst,matrix_A[8868],matrix_B[68],mul_res1[8868]);
multi_7x28 multi_7x28_mod_8869(clk,rst,matrix_A[8869],matrix_B[69],mul_res1[8869]);
multi_7x28 multi_7x28_mod_8870(clk,rst,matrix_A[8870],matrix_B[70],mul_res1[8870]);
multi_7x28 multi_7x28_mod_8871(clk,rst,matrix_A[8871],matrix_B[71],mul_res1[8871]);
multi_7x28 multi_7x28_mod_8872(clk,rst,matrix_A[8872],matrix_B[72],mul_res1[8872]);
multi_7x28 multi_7x28_mod_8873(clk,rst,matrix_A[8873],matrix_B[73],mul_res1[8873]);
multi_7x28 multi_7x28_mod_8874(clk,rst,matrix_A[8874],matrix_B[74],mul_res1[8874]);
multi_7x28 multi_7x28_mod_8875(clk,rst,matrix_A[8875],matrix_B[75],mul_res1[8875]);
multi_7x28 multi_7x28_mod_8876(clk,rst,matrix_A[8876],matrix_B[76],mul_res1[8876]);
multi_7x28 multi_7x28_mod_8877(clk,rst,matrix_A[8877],matrix_B[77],mul_res1[8877]);
multi_7x28 multi_7x28_mod_8878(clk,rst,matrix_A[8878],matrix_B[78],mul_res1[8878]);
multi_7x28 multi_7x28_mod_8879(clk,rst,matrix_A[8879],matrix_B[79],mul_res1[8879]);
multi_7x28 multi_7x28_mod_8880(clk,rst,matrix_A[8880],matrix_B[80],mul_res1[8880]);
multi_7x28 multi_7x28_mod_8881(clk,rst,matrix_A[8881],matrix_B[81],mul_res1[8881]);
multi_7x28 multi_7x28_mod_8882(clk,rst,matrix_A[8882],matrix_B[82],mul_res1[8882]);
multi_7x28 multi_7x28_mod_8883(clk,rst,matrix_A[8883],matrix_B[83],mul_res1[8883]);
multi_7x28 multi_7x28_mod_8884(clk,rst,matrix_A[8884],matrix_B[84],mul_res1[8884]);
multi_7x28 multi_7x28_mod_8885(clk,rst,matrix_A[8885],matrix_B[85],mul_res1[8885]);
multi_7x28 multi_7x28_mod_8886(clk,rst,matrix_A[8886],matrix_B[86],mul_res1[8886]);
multi_7x28 multi_7x28_mod_8887(clk,rst,matrix_A[8887],matrix_B[87],mul_res1[8887]);
multi_7x28 multi_7x28_mod_8888(clk,rst,matrix_A[8888],matrix_B[88],mul_res1[8888]);
multi_7x28 multi_7x28_mod_8889(clk,rst,matrix_A[8889],matrix_B[89],mul_res1[8889]);
multi_7x28 multi_7x28_mod_8890(clk,rst,matrix_A[8890],matrix_B[90],mul_res1[8890]);
multi_7x28 multi_7x28_mod_8891(clk,rst,matrix_A[8891],matrix_B[91],mul_res1[8891]);
multi_7x28 multi_7x28_mod_8892(clk,rst,matrix_A[8892],matrix_B[92],mul_res1[8892]);
multi_7x28 multi_7x28_mod_8893(clk,rst,matrix_A[8893],matrix_B[93],mul_res1[8893]);
multi_7x28 multi_7x28_mod_8894(clk,rst,matrix_A[8894],matrix_B[94],mul_res1[8894]);
multi_7x28 multi_7x28_mod_8895(clk,rst,matrix_A[8895],matrix_B[95],mul_res1[8895]);
multi_7x28 multi_7x28_mod_8896(clk,rst,matrix_A[8896],matrix_B[96],mul_res1[8896]);
multi_7x28 multi_7x28_mod_8897(clk,rst,matrix_A[8897],matrix_B[97],mul_res1[8897]);
multi_7x28 multi_7x28_mod_8898(clk,rst,matrix_A[8898],matrix_B[98],mul_res1[8898]);
multi_7x28 multi_7x28_mod_8899(clk,rst,matrix_A[8899],matrix_B[99],mul_res1[8899]);
multi_7x28 multi_7x28_mod_8900(clk,rst,matrix_A[8900],matrix_B[100],mul_res1[8900]);
multi_7x28 multi_7x28_mod_8901(clk,rst,matrix_A[8901],matrix_B[101],mul_res1[8901]);
multi_7x28 multi_7x28_mod_8902(clk,rst,matrix_A[8902],matrix_B[102],mul_res1[8902]);
multi_7x28 multi_7x28_mod_8903(clk,rst,matrix_A[8903],matrix_B[103],mul_res1[8903]);
multi_7x28 multi_7x28_mod_8904(clk,rst,matrix_A[8904],matrix_B[104],mul_res1[8904]);
multi_7x28 multi_7x28_mod_8905(clk,rst,matrix_A[8905],matrix_B[105],mul_res1[8905]);
multi_7x28 multi_7x28_mod_8906(clk,rst,matrix_A[8906],matrix_B[106],mul_res1[8906]);
multi_7x28 multi_7x28_mod_8907(clk,rst,matrix_A[8907],matrix_B[107],mul_res1[8907]);
multi_7x28 multi_7x28_mod_8908(clk,rst,matrix_A[8908],matrix_B[108],mul_res1[8908]);
multi_7x28 multi_7x28_mod_8909(clk,rst,matrix_A[8909],matrix_B[109],mul_res1[8909]);
multi_7x28 multi_7x28_mod_8910(clk,rst,matrix_A[8910],matrix_B[110],mul_res1[8910]);
multi_7x28 multi_7x28_mod_8911(clk,rst,matrix_A[8911],matrix_B[111],mul_res1[8911]);
multi_7x28 multi_7x28_mod_8912(clk,rst,matrix_A[8912],matrix_B[112],mul_res1[8912]);
multi_7x28 multi_7x28_mod_8913(clk,rst,matrix_A[8913],matrix_B[113],mul_res1[8913]);
multi_7x28 multi_7x28_mod_8914(clk,rst,matrix_A[8914],matrix_B[114],mul_res1[8914]);
multi_7x28 multi_7x28_mod_8915(clk,rst,matrix_A[8915],matrix_B[115],mul_res1[8915]);
multi_7x28 multi_7x28_mod_8916(clk,rst,matrix_A[8916],matrix_B[116],mul_res1[8916]);
multi_7x28 multi_7x28_mod_8917(clk,rst,matrix_A[8917],matrix_B[117],mul_res1[8917]);
multi_7x28 multi_7x28_mod_8918(clk,rst,matrix_A[8918],matrix_B[118],mul_res1[8918]);
multi_7x28 multi_7x28_mod_8919(clk,rst,matrix_A[8919],matrix_B[119],mul_res1[8919]);
multi_7x28 multi_7x28_mod_8920(clk,rst,matrix_A[8920],matrix_B[120],mul_res1[8920]);
multi_7x28 multi_7x28_mod_8921(clk,rst,matrix_A[8921],matrix_B[121],mul_res1[8921]);
multi_7x28 multi_7x28_mod_8922(clk,rst,matrix_A[8922],matrix_B[122],mul_res1[8922]);
multi_7x28 multi_7x28_mod_8923(clk,rst,matrix_A[8923],matrix_B[123],mul_res1[8923]);
multi_7x28 multi_7x28_mod_8924(clk,rst,matrix_A[8924],matrix_B[124],mul_res1[8924]);
multi_7x28 multi_7x28_mod_8925(clk,rst,matrix_A[8925],matrix_B[125],mul_res1[8925]);
multi_7x28 multi_7x28_mod_8926(clk,rst,matrix_A[8926],matrix_B[126],mul_res1[8926]);
multi_7x28 multi_7x28_mod_8927(clk,rst,matrix_A[8927],matrix_B[127],mul_res1[8927]);
multi_7x28 multi_7x28_mod_8928(clk,rst,matrix_A[8928],matrix_B[128],mul_res1[8928]);
multi_7x28 multi_7x28_mod_8929(clk,rst,matrix_A[8929],matrix_B[129],mul_res1[8929]);
multi_7x28 multi_7x28_mod_8930(clk,rst,matrix_A[8930],matrix_B[130],mul_res1[8930]);
multi_7x28 multi_7x28_mod_8931(clk,rst,matrix_A[8931],matrix_B[131],mul_res1[8931]);
multi_7x28 multi_7x28_mod_8932(clk,rst,matrix_A[8932],matrix_B[132],mul_res1[8932]);
multi_7x28 multi_7x28_mod_8933(clk,rst,matrix_A[8933],matrix_B[133],mul_res1[8933]);
multi_7x28 multi_7x28_mod_8934(clk,rst,matrix_A[8934],matrix_B[134],mul_res1[8934]);
multi_7x28 multi_7x28_mod_8935(clk,rst,matrix_A[8935],matrix_B[135],mul_res1[8935]);
multi_7x28 multi_7x28_mod_8936(clk,rst,matrix_A[8936],matrix_B[136],mul_res1[8936]);
multi_7x28 multi_7x28_mod_8937(clk,rst,matrix_A[8937],matrix_B[137],mul_res1[8937]);
multi_7x28 multi_7x28_mod_8938(clk,rst,matrix_A[8938],matrix_B[138],mul_res1[8938]);
multi_7x28 multi_7x28_mod_8939(clk,rst,matrix_A[8939],matrix_B[139],mul_res1[8939]);
multi_7x28 multi_7x28_mod_8940(clk,rst,matrix_A[8940],matrix_B[140],mul_res1[8940]);
multi_7x28 multi_7x28_mod_8941(clk,rst,matrix_A[8941],matrix_B[141],mul_res1[8941]);
multi_7x28 multi_7x28_mod_8942(clk,rst,matrix_A[8942],matrix_B[142],mul_res1[8942]);
multi_7x28 multi_7x28_mod_8943(clk,rst,matrix_A[8943],matrix_B[143],mul_res1[8943]);
multi_7x28 multi_7x28_mod_8944(clk,rst,matrix_A[8944],matrix_B[144],mul_res1[8944]);
multi_7x28 multi_7x28_mod_8945(clk,rst,matrix_A[8945],matrix_B[145],mul_res1[8945]);
multi_7x28 multi_7x28_mod_8946(clk,rst,matrix_A[8946],matrix_B[146],mul_res1[8946]);
multi_7x28 multi_7x28_mod_8947(clk,rst,matrix_A[8947],matrix_B[147],mul_res1[8947]);
multi_7x28 multi_7x28_mod_8948(clk,rst,matrix_A[8948],matrix_B[148],mul_res1[8948]);
multi_7x28 multi_7x28_mod_8949(clk,rst,matrix_A[8949],matrix_B[149],mul_res1[8949]);
multi_7x28 multi_7x28_mod_8950(clk,rst,matrix_A[8950],matrix_B[150],mul_res1[8950]);
multi_7x28 multi_7x28_mod_8951(clk,rst,matrix_A[8951],matrix_B[151],mul_res1[8951]);
multi_7x28 multi_7x28_mod_8952(clk,rst,matrix_A[8952],matrix_B[152],mul_res1[8952]);
multi_7x28 multi_7x28_mod_8953(clk,rst,matrix_A[8953],matrix_B[153],mul_res1[8953]);
multi_7x28 multi_7x28_mod_8954(clk,rst,matrix_A[8954],matrix_B[154],mul_res1[8954]);
multi_7x28 multi_7x28_mod_8955(clk,rst,matrix_A[8955],matrix_B[155],mul_res1[8955]);
multi_7x28 multi_7x28_mod_8956(clk,rst,matrix_A[8956],matrix_B[156],mul_res1[8956]);
multi_7x28 multi_7x28_mod_8957(clk,rst,matrix_A[8957],matrix_B[157],mul_res1[8957]);
multi_7x28 multi_7x28_mod_8958(clk,rst,matrix_A[8958],matrix_B[158],mul_res1[8958]);
multi_7x28 multi_7x28_mod_8959(clk,rst,matrix_A[8959],matrix_B[159],mul_res1[8959]);
multi_7x28 multi_7x28_mod_8960(clk,rst,matrix_A[8960],matrix_B[160],mul_res1[8960]);
multi_7x28 multi_7x28_mod_8961(clk,rst,matrix_A[8961],matrix_B[161],mul_res1[8961]);
multi_7x28 multi_7x28_mod_8962(clk,rst,matrix_A[8962],matrix_B[162],mul_res1[8962]);
multi_7x28 multi_7x28_mod_8963(clk,rst,matrix_A[8963],matrix_B[163],mul_res1[8963]);
multi_7x28 multi_7x28_mod_8964(clk,rst,matrix_A[8964],matrix_B[164],mul_res1[8964]);
multi_7x28 multi_7x28_mod_8965(clk,rst,matrix_A[8965],matrix_B[165],mul_res1[8965]);
multi_7x28 multi_7x28_mod_8966(clk,rst,matrix_A[8966],matrix_B[166],mul_res1[8966]);
multi_7x28 multi_7x28_mod_8967(clk,rst,matrix_A[8967],matrix_B[167],mul_res1[8967]);
multi_7x28 multi_7x28_mod_8968(clk,rst,matrix_A[8968],matrix_B[168],mul_res1[8968]);
multi_7x28 multi_7x28_mod_8969(clk,rst,matrix_A[8969],matrix_B[169],mul_res1[8969]);
multi_7x28 multi_7x28_mod_8970(clk,rst,matrix_A[8970],matrix_B[170],mul_res1[8970]);
multi_7x28 multi_7x28_mod_8971(clk,rst,matrix_A[8971],matrix_B[171],mul_res1[8971]);
multi_7x28 multi_7x28_mod_8972(clk,rst,matrix_A[8972],matrix_B[172],mul_res1[8972]);
multi_7x28 multi_7x28_mod_8973(clk,rst,matrix_A[8973],matrix_B[173],mul_res1[8973]);
multi_7x28 multi_7x28_mod_8974(clk,rst,matrix_A[8974],matrix_B[174],mul_res1[8974]);
multi_7x28 multi_7x28_mod_8975(clk,rst,matrix_A[8975],matrix_B[175],mul_res1[8975]);
multi_7x28 multi_7x28_mod_8976(clk,rst,matrix_A[8976],matrix_B[176],mul_res1[8976]);
multi_7x28 multi_7x28_mod_8977(clk,rst,matrix_A[8977],matrix_B[177],mul_res1[8977]);
multi_7x28 multi_7x28_mod_8978(clk,rst,matrix_A[8978],matrix_B[178],mul_res1[8978]);
multi_7x28 multi_7x28_mod_8979(clk,rst,matrix_A[8979],matrix_B[179],mul_res1[8979]);
multi_7x28 multi_7x28_mod_8980(clk,rst,matrix_A[8980],matrix_B[180],mul_res1[8980]);
multi_7x28 multi_7x28_mod_8981(clk,rst,matrix_A[8981],matrix_B[181],mul_res1[8981]);
multi_7x28 multi_7x28_mod_8982(clk,rst,matrix_A[8982],matrix_B[182],mul_res1[8982]);
multi_7x28 multi_7x28_mod_8983(clk,rst,matrix_A[8983],matrix_B[183],mul_res1[8983]);
multi_7x28 multi_7x28_mod_8984(clk,rst,matrix_A[8984],matrix_B[184],mul_res1[8984]);
multi_7x28 multi_7x28_mod_8985(clk,rst,matrix_A[8985],matrix_B[185],mul_res1[8985]);
multi_7x28 multi_7x28_mod_8986(clk,rst,matrix_A[8986],matrix_B[186],mul_res1[8986]);
multi_7x28 multi_7x28_mod_8987(clk,rst,matrix_A[8987],matrix_B[187],mul_res1[8987]);
multi_7x28 multi_7x28_mod_8988(clk,rst,matrix_A[8988],matrix_B[188],mul_res1[8988]);
multi_7x28 multi_7x28_mod_8989(clk,rst,matrix_A[8989],matrix_B[189],mul_res1[8989]);
multi_7x28 multi_7x28_mod_8990(clk,rst,matrix_A[8990],matrix_B[190],mul_res1[8990]);
multi_7x28 multi_7x28_mod_8991(clk,rst,matrix_A[8991],matrix_B[191],mul_res1[8991]);
multi_7x28 multi_7x28_mod_8992(clk,rst,matrix_A[8992],matrix_B[192],mul_res1[8992]);
multi_7x28 multi_7x28_mod_8993(clk,rst,matrix_A[8993],matrix_B[193],mul_res1[8993]);
multi_7x28 multi_7x28_mod_8994(clk,rst,matrix_A[8994],matrix_B[194],mul_res1[8994]);
multi_7x28 multi_7x28_mod_8995(clk,rst,matrix_A[8995],matrix_B[195],mul_res1[8995]);
multi_7x28 multi_7x28_mod_8996(clk,rst,matrix_A[8996],matrix_B[196],mul_res1[8996]);
multi_7x28 multi_7x28_mod_8997(clk,rst,matrix_A[8997],matrix_B[197],mul_res1[8997]);
multi_7x28 multi_7x28_mod_8998(clk,rst,matrix_A[8998],matrix_B[198],mul_res1[8998]);
multi_7x28 multi_7x28_mod_8999(clk,rst,matrix_A[8999],matrix_B[199],mul_res1[8999]);
multi_7x28 multi_7x28_mod_9000(clk,rst,matrix_A[9000],matrix_B[0],mul_res1[9000]);
multi_7x28 multi_7x28_mod_9001(clk,rst,matrix_A[9001],matrix_B[1],mul_res1[9001]);
multi_7x28 multi_7x28_mod_9002(clk,rst,matrix_A[9002],matrix_B[2],mul_res1[9002]);
multi_7x28 multi_7x28_mod_9003(clk,rst,matrix_A[9003],matrix_B[3],mul_res1[9003]);
multi_7x28 multi_7x28_mod_9004(clk,rst,matrix_A[9004],matrix_B[4],mul_res1[9004]);
multi_7x28 multi_7x28_mod_9005(clk,rst,matrix_A[9005],matrix_B[5],mul_res1[9005]);
multi_7x28 multi_7x28_mod_9006(clk,rst,matrix_A[9006],matrix_B[6],mul_res1[9006]);
multi_7x28 multi_7x28_mod_9007(clk,rst,matrix_A[9007],matrix_B[7],mul_res1[9007]);
multi_7x28 multi_7x28_mod_9008(clk,rst,matrix_A[9008],matrix_B[8],mul_res1[9008]);
multi_7x28 multi_7x28_mod_9009(clk,rst,matrix_A[9009],matrix_B[9],mul_res1[9009]);
multi_7x28 multi_7x28_mod_9010(clk,rst,matrix_A[9010],matrix_B[10],mul_res1[9010]);
multi_7x28 multi_7x28_mod_9011(clk,rst,matrix_A[9011],matrix_B[11],mul_res1[9011]);
multi_7x28 multi_7x28_mod_9012(clk,rst,matrix_A[9012],matrix_B[12],mul_res1[9012]);
multi_7x28 multi_7x28_mod_9013(clk,rst,matrix_A[9013],matrix_B[13],mul_res1[9013]);
multi_7x28 multi_7x28_mod_9014(clk,rst,matrix_A[9014],matrix_B[14],mul_res1[9014]);
multi_7x28 multi_7x28_mod_9015(clk,rst,matrix_A[9015],matrix_B[15],mul_res1[9015]);
multi_7x28 multi_7x28_mod_9016(clk,rst,matrix_A[9016],matrix_B[16],mul_res1[9016]);
multi_7x28 multi_7x28_mod_9017(clk,rst,matrix_A[9017],matrix_B[17],mul_res1[9017]);
multi_7x28 multi_7x28_mod_9018(clk,rst,matrix_A[9018],matrix_B[18],mul_res1[9018]);
multi_7x28 multi_7x28_mod_9019(clk,rst,matrix_A[9019],matrix_B[19],mul_res1[9019]);
multi_7x28 multi_7x28_mod_9020(clk,rst,matrix_A[9020],matrix_B[20],mul_res1[9020]);
multi_7x28 multi_7x28_mod_9021(clk,rst,matrix_A[9021],matrix_B[21],mul_res1[9021]);
multi_7x28 multi_7x28_mod_9022(clk,rst,matrix_A[9022],matrix_B[22],mul_res1[9022]);
multi_7x28 multi_7x28_mod_9023(clk,rst,matrix_A[9023],matrix_B[23],mul_res1[9023]);
multi_7x28 multi_7x28_mod_9024(clk,rst,matrix_A[9024],matrix_B[24],mul_res1[9024]);
multi_7x28 multi_7x28_mod_9025(clk,rst,matrix_A[9025],matrix_B[25],mul_res1[9025]);
multi_7x28 multi_7x28_mod_9026(clk,rst,matrix_A[9026],matrix_B[26],mul_res1[9026]);
multi_7x28 multi_7x28_mod_9027(clk,rst,matrix_A[9027],matrix_B[27],mul_res1[9027]);
multi_7x28 multi_7x28_mod_9028(clk,rst,matrix_A[9028],matrix_B[28],mul_res1[9028]);
multi_7x28 multi_7x28_mod_9029(clk,rst,matrix_A[9029],matrix_B[29],mul_res1[9029]);
multi_7x28 multi_7x28_mod_9030(clk,rst,matrix_A[9030],matrix_B[30],mul_res1[9030]);
multi_7x28 multi_7x28_mod_9031(clk,rst,matrix_A[9031],matrix_B[31],mul_res1[9031]);
multi_7x28 multi_7x28_mod_9032(clk,rst,matrix_A[9032],matrix_B[32],mul_res1[9032]);
multi_7x28 multi_7x28_mod_9033(clk,rst,matrix_A[9033],matrix_B[33],mul_res1[9033]);
multi_7x28 multi_7x28_mod_9034(clk,rst,matrix_A[9034],matrix_B[34],mul_res1[9034]);
multi_7x28 multi_7x28_mod_9035(clk,rst,matrix_A[9035],matrix_B[35],mul_res1[9035]);
multi_7x28 multi_7x28_mod_9036(clk,rst,matrix_A[9036],matrix_B[36],mul_res1[9036]);
multi_7x28 multi_7x28_mod_9037(clk,rst,matrix_A[9037],matrix_B[37],mul_res1[9037]);
multi_7x28 multi_7x28_mod_9038(clk,rst,matrix_A[9038],matrix_B[38],mul_res1[9038]);
multi_7x28 multi_7x28_mod_9039(clk,rst,matrix_A[9039],matrix_B[39],mul_res1[9039]);
multi_7x28 multi_7x28_mod_9040(clk,rst,matrix_A[9040],matrix_B[40],mul_res1[9040]);
multi_7x28 multi_7x28_mod_9041(clk,rst,matrix_A[9041],matrix_B[41],mul_res1[9041]);
multi_7x28 multi_7x28_mod_9042(clk,rst,matrix_A[9042],matrix_B[42],mul_res1[9042]);
multi_7x28 multi_7x28_mod_9043(clk,rst,matrix_A[9043],matrix_B[43],mul_res1[9043]);
multi_7x28 multi_7x28_mod_9044(clk,rst,matrix_A[9044],matrix_B[44],mul_res1[9044]);
multi_7x28 multi_7x28_mod_9045(clk,rst,matrix_A[9045],matrix_B[45],mul_res1[9045]);
multi_7x28 multi_7x28_mod_9046(clk,rst,matrix_A[9046],matrix_B[46],mul_res1[9046]);
multi_7x28 multi_7x28_mod_9047(clk,rst,matrix_A[9047],matrix_B[47],mul_res1[9047]);
multi_7x28 multi_7x28_mod_9048(clk,rst,matrix_A[9048],matrix_B[48],mul_res1[9048]);
multi_7x28 multi_7x28_mod_9049(clk,rst,matrix_A[9049],matrix_B[49],mul_res1[9049]);
multi_7x28 multi_7x28_mod_9050(clk,rst,matrix_A[9050],matrix_B[50],mul_res1[9050]);
multi_7x28 multi_7x28_mod_9051(clk,rst,matrix_A[9051],matrix_B[51],mul_res1[9051]);
multi_7x28 multi_7x28_mod_9052(clk,rst,matrix_A[9052],matrix_B[52],mul_res1[9052]);
multi_7x28 multi_7x28_mod_9053(clk,rst,matrix_A[9053],matrix_B[53],mul_res1[9053]);
multi_7x28 multi_7x28_mod_9054(clk,rst,matrix_A[9054],matrix_B[54],mul_res1[9054]);
multi_7x28 multi_7x28_mod_9055(clk,rst,matrix_A[9055],matrix_B[55],mul_res1[9055]);
multi_7x28 multi_7x28_mod_9056(clk,rst,matrix_A[9056],matrix_B[56],mul_res1[9056]);
multi_7x28 multi_7x28_mod_9057(clk,rst,matrix_A[9057],matrix_B[57],mul_res1[9057]);
multi_7x28 multi_7x28_mod_9058(clk,rst,matrix_A[9058],matrix_B[58],mul_res1[9058]);
multi_7x28 multi_7x28_mod_9059(clk,rst,matrix_A[9059],matrix_B[59],mul_res1[9059]);
multi_7x28 multi_7x28_mod_9060(clk,rst,matrix_A[9060],matrix_B[60],mul_res1[9060]);
multi_7x28 multi_7x28_mod_9061(clk,rst,matrix_A[9061],matrix_B[61],mul_res1[9061]);
multi_7x28 multi_7x28_mod_9062(clk,rst,matrix_A[9062],matrix_B[62],mul_res1[9062]);
multi_7x28 multi_7x28_mod_9063(clk,rst,matrix_A[9063],matrix_B[63],mul_res1[9063]);
multi_7x28 multi_7x28_mod_9064(clk,rst,matrix_A[9064],matrix_B[64],mul_res1[9064]);
multi_7x28 multi_7x28_mod_9065(clk,rst,matrix_A[9065],matrix_B[65],mul_res1[9065]);
multi_7x28 multi_7x28_mod_9066(clk,rst,matrix_A[9066],matrix_B[66],mul_res1[9066]);
multi_7x28 multi_7x28_mod_9067(clk,rst,matrix_A[9067],matrix_B[67],mul_res1[9067]);
multi_7x28 multi_7x28_mod_9068(clk,rst,matrix_A[9068],matrix_B[68],mul_res1[9068]);
multi_7x28 multi_7x28_mod_9069(clk,rst,matrix_A[9069],matrix_B[69],mul_res1[9069]);
multi_7x28 multi_7x28_mod_9070(clk,rst,matrix_A[9070],matrix_B[70],mul_res1[9070]);
multi_7x28 multi_7x28_mod_9071(clk,rst,matrix_A[9071],matrix_B[71],mul_res1[9071]);
multi_7x28 multi_7x28_mod_9072(clk,rst,matrix_A[9072],matrix_B[72],mul_res1[9072]);
multi_7x28 multi_7x28_mod_9073(clk,rst,matrix_A[9073],matrix_B[73],mul_res1[9073]);
multi_7x28 multi_7x28_mod_9074(clk,rst,matrix_A[9074],matrix_B[74],mul_res1[9074]);
multi_7x28 multi_7x28_mod_9075(clk,rst,matrix_A[9075],matrix_B[75],mul_res1[9075]);
multi_7x28 multi_7x28_mod_9076(clk,rst,matrix_A[9076],matrix_B[76],mul_res1[9076]);
multi_7x28 multi_7x28_mod_9077(clk,rst,matrix_A[9077],matrix_B[77],mul_res1[9077]);
multi_7x28 multi_7x28_mod_9078(clk,rst,matrix_A[9078],matrix_B[78],mul_res1[9078]);
multi_7x28 multi_7x28_mod_9079(clk,rst,matrix_A[9079],matrix_B[79],mul_res1[9079]);
multi_7x28 multi_7x28_mod_9080(clk,rst,matrix_A[9080],matrix_B[80],mul_res1[9080]);
multi_7x28 multi_7x28_mod_9081(clk,rst,matrix_A[9081],matrix_B[81],mul_res1[9081]);
multi_7x28 multi_7x28_mod_9082(clk,rst,matrix_A[9082],matrix_B[82],mul_res1[9082]);
multi_7x28 multi_7x28_mod_9083(clk,rst,matrix_A[9083],matrix_B[83],mul_res1[9083]);
multi_7x28 multi_7x28_mod_9084(clk,rst,matrix_A[9084],matrix_B[84],mul_res1[9084]);
multi_7x28 multi_7x28_mod_9085(clk,rst,matrix_A[9085],matrix_B[85],mul_res1[9085]);
multi_7x28 multi_7x28_mod_9086(clk,rst,matrix_A[9086],matrix_B[86],mul_res1[9086]);
multi_7x28 multi_7x28_mod_9087(clk,rst,matrix_A[9087],matrix_B[87],mul_res1[9087]);
multi_7x28 multi_7x28_mod_9088(clk,rst,matrix_A[9088],matrix_B[88],mul_res1[9088]);
multi_7x28 multi_7x28_mod_9089(clk,rst,matrix_A[9089],matrix_B[89],mul_res1[9089]);
multi_7x28 multi_7x28_mod_9090(clk,rst,matrix_A[9090],matrix_B[90],mul_res1[9090]);
multi_7x28 multi_7x28_mod_9091(clk,rst,matrix_A[9091],matrix_B[91],mul_res1[9091]);
multi_7x28 multi_7x28_mod_9092(clk,rst,matrix_A[9092],matrix_B[92],mul_res1[9092]);
multi_7x28 multi_7x28_mod_9093(clk,rst,matrix_A[9093],matrix_B[93],mul_res1[9093]);
multi_7x28 multi_7x28_mod_9094(clk,rst,matrix_A[9094],matrix_B[94],mul_res1[9094]);
multi_7x28 multi_7x28_mod_9095(clk,rst,matrix_A[9095],matrix_B[95],mul_res1[9095]);
multi_7x28 multi_7x28_mod_9096(clk,rst,matrix_A[9096],matrix_B[96],mul_res1[9096]);
multi_7x28 multi_7x28_mod_9097(clk,rst,matrix_A[9097],matrix_B[97],mul_res1[9097]);
multi_7x28 multi_7x28_mod_9098(clk,rst,matrix_A[9098],matrix_B[98],mul_res1[9098]);
multi_7x28 multi_7x28_mod_9099(clk,rst,matrix_A[9099],matrix_B[99],mul_res1[9099]);
multi_7x28 multi_7x28_mod_9100(clk,rst,matrix_A[9100],matrix_B[100],mul_res1[9100]);
multi_7x28 multi_7x28_mod_9101(clk,rst,matrix_A[9101],matrix_B[101],mul_res1[9101]);
multi_7x28 multi_7x28_mod_9102(clk,rst,matrix_A[9102],matrix_B[102],mul_res1[9102]);
multi_7x28 multi_7x28_mod_9103(clk,rst,matrix_A[9103],matrix_B[103],mul_res1[9103]);
multi_7x28 multi_7x28_mod_9104(clk,rst,matrix_A[9104],matrix_B[104],mul_res1[9104]);
multi_7x28 multi_7x28_mod_9105(clk,rst,matrix_A[9105],matrix_B[105],mul_res1[9105]);
multi_7x28 multi_7x28_mod_9106(clk,rst,matrix_A[9106],matrix_B[106],mul_res1[9106]);
multi_7x28 multi_7x28_mod_9107(clk,rst,matrix_A[9107],matrix_B[107],mul_res1[9107]);
multi_7x28 multi_7x28_mod_9108(clk,rst,matrix_A[9108],matrix_B[108],mul_res1[9108]);
multi_7x28 multi_7x28_mod_9109(clk,rst,matrix_A[9109],matrix_B[109],mul_res1[9109]);
multi_7x28 multi_7x28_mod_9110(clk,rst,matrix_A[9110],matrix_B[110],mul_res1[9110]);
multi_7x28 multi_7x28_mod_9111(clk,rst,matrix_A[9111],matrix_B[111],mul_res1[9111]);
multi_7x28 multi_7x28_mod_9112(clk,rst,matrix_A[9112],matrix_B[112],mul_res1[9112]);
multi_7x28 multi_7x28_mod_9113(clk,rst,matrix_A[9113],matrix_B[113],mul_res1[9113]);
multi_7x28 multi_7x28_mod_9114(clk,rst,matrix_A[9114],matrix_B[114],mul_res1[9114]);
multi_7x28 multi_7x28_mod_9115(clk,rst,matrix_A[9115],matrix_B[115],mul_res1[9115]);
multi_7x28 multi_7x28_mod_9116(clk,rst,matrix_A[9116],matrix_B[116],mul_res1[9116]);
multi_7x28 multi_7x28_mod_9117(clk,rst,matrix_A[9117],matrix_B[117],mul_res1[9117]);
multi_7x28 multi_7x28_mod_9118(clk,rst,matrix_A[9118],matrix_B[118],mul_res1[9118]);
multi_7x28 multi_7x28_mod_9119(clk,rst,matrix_A[9119],matrix_B[119],mul_res1[9119]);
multi_7x28 multi_7x28_mod_9120(clk,rst,matrix_A[9120],matrix_B[120],mul_res1[9120]);
multi_7x28 multi_7x28_mod_9121(clk,rst,matrix_A[9121],matrix_B[121],mul_res1[9121]);
multi_7x28 multi_7x28_mod_9122(clk,rst,matrix_A[9122],matrix_B[122],mul_res1[9122]);
multi_7x28 multi_7x28_mod_9123(clk,rst,matrix_A[9123],matrix_B[123],mul_res1[9123]);
multi_7x28 multi_7x28_mod_9124(clk,rst,matrix_A[9124],matrix_B[124],mul_res1[9124]);
multi_7x28 multi_7x28_mod_9125(clk,rst,matrix_A[9125],matrix_B[125],mul_res1[9125]);
multi_7x28 multi_7x28_mod_9126(clk,rst,matrix_A[9126],matrix_B[126],mul_res1[9126]);
multi_7x28 multi_7x28_mod_9127(clk,rst,matrix_A[9127],matrix_B[127],mul_res1[9127]);
multi_7x28 multi_7x28_mod_9128(clk,rst,matrix_A[9128],matrix_B[128],mul_res1[9128]);
multi_7x28 multi_7x28_mod_9129(clk,rst,matrix_A[9129],matrix_B[129],mul_res1[9129]);
multi_7x28 multi_7x28_mod_9130(clk,rst,matrix_A[9130],matrix_B[130],mul_res1[9130]);
multi_7x28 multi_7x28_mod_9131(clk,rst,matrix_A[9131],matrix_B[131],mul_res1[9131]);
multi_7x28 multi_7x28_mod_9132(clk,rst,matrix_A[9132],matrix_B[132],mul_res1[9132]);
multi_7x28 multi_7x28_mod_9133(clk,rst,matrix_A[9133],matrix_B[133],mul_res1[9133]);
multi_7x28 multi_7x28_mod_9134(clk,rst,matrix_A[9134],matrix_B[134],mul_res1[9134]);
multi_7x28 multi_7x28_mod_9135(clk,rst,matrix_A[9135],matrix_B[135],mul_res1[9135]);
multi_7x28 multi_7x28_mod_9136(clk,rst,matrix_A[9136],matrix_B[136],mul_res1[9136]);
multi_7x28 multi_7x28_mod_9137(clk,rst,matrix_A[9137],matrix_B[137],mul_res1[9137]);
multi_7x28 multi_7x28_mod_9138(clk,rst,matrix_A[9138],matrix_B[138],mul_res1[9138]);
multi_7x28 multi_7x28_mod_9139(clk,rst,matrix_A[9139],matrix_B[139],mul_res1[9139]);
multi_7x28 multi_7x28_mod_9140(clk,rst,matrix_A[9140],matrix_B[140],mul_res1[9140]);
multi_7x28 multi_7x28_mod_9141(clk,rst,matrix_A[9141],matrix_B[141],mul_res1[9141]);
multi_7x28 multi_7x28_mod_9142(clk,rst,matrix_A[9142],matrix_B[142],mul_res1[9142]);
multi_7x28 multi_7x28_mod_9143(clk,rst,matrix_A[9143],matrix_B[143],mul_res1[9143]);
multi_7x28 multi_7x28_mod_9144(clk,rst,matrix_A[9144],matrix_B[144],mul_res1[9144]);
multi_7x28 multi_7x28_mod_9145(clk,rst,matrix_A[9145],matrix_B[145],mul_res1[9145]);
multi_7x28 multi_7x28_mod_9146(clk,rst,matrix_A[9146],matrix_B[146],mul_res1[9146]);
multi_7x28 multi_7x28_mod_9147(clk,rst,matrix_A[9147],matrix_B[147],mul_res1[9147]);
multi_7x28 multi_7x28_mod_9148(clk,rst,matrix_A[9148],matrix_B[148],mul_res1[9148]);
multi_7x28 multi_7x28_mod_9149(clk,rst,matrix_A[9149],matrix_B[149],mul_res1[9149]);
multi_7x28 multi_7x28_mod_9150(clk,rst,matrix_A[9150],matrix_B[150],mul_res1[9150]);
multi_7x28 multi_7x28_mod_9151(clk,rst,matrix_A[9151],matrix_B[151],mul_res1[9151]);
multi_7x28 multi_7x28_mod_9152(clk,rst,matrix_A[9152],matrix_B[152],mul_res1[9152]);
multi_7x28 multi_7x28_mod_9153(clk,rst,matrix_A[9153],matrix_B[153],mul_res1[9153]);
multi_7x28 multi_7x28_mod_9154(clk,rst,matrix_A[9154],matrix_B[154],mul_res1[9154]);
multi_7x28 multi_7x28_mod_9155(clk,rst,matrix_A[9155],matrix_B[155],mul_res1[9155]);
multi_7x28 multi_7x28_mod_9156(clk,rst,matrix_A[9156],matrix_B[156],mul_res1[9156]);
multi_7x28 multi_7x28_mod_9157(clk,rst,matrix_A[9157],matrix_B[157],mul_res1[9157]);
multi_7x28 multi_7x28_mod_9158(clk,rst,matrix_A[9158],matrix_B[158],mul_res1[9158]);
multi_7x28 multi_7x28_mod_9159(clk,rst,matrix_A[9159],matrix_B[159],mul_res1[9159]);
multi_7x28 multi_7x28_mod_9160(clk,rst,matrix_A[9160],matrix_B[160],mul_res1[9160]);
multi_7x28 multi_7x28_mod_9161(clk,rst,matrix_A[9161],matrix_B[161],mul_res1[9161]);
multi_7x28 multi_7x28_mod_9162(clk,rst,matrix_A[9162],matrix_B[162],mul_res1[9162]);
multi_7x28 multi_7x28_mod_9163(clk,rst,matrix_A[9163],matrix_B[163],mul_res1[9163]);
multi_7x28 multi_7x28_mod_9164(clk,rst,matrix_A[9164],matrix_B[164],mul_res1[9164]);
multi_7x28 multi_7x28_mod_9165(clk,rst,matrix_A[9165],matrix_B[165],mul_res1[9165]);
multi_7x28 multi_7x28_mod_9166(clk,rst,matrix_A[9166],matrix_B[166],mul_res1[9166]);
multi_7x28 multi_7x28_mod_9167(clk,rst,matrix_A[9167],matrix_B[167],mul_res1[9167]);
multi_7x28 multi_7x28_mod_9168(clk,rst,matrix_A[9168],matrix_B[168],mul_res1[9168]);
multi_7x28 multi_7x28_mod_9169(clk,rst,matrix_A[9169],matrix_B[169],mul_res1[9169]);
multi_7x28 multi_7x28_mod_9170(clk,rst,matrix_A[9170],matrix_B[170],mul_res1[9170]);
multi_7x28 multi_7x28_mod_9171(clk,rst,matrix_A[9171],matrix_B[171],mul_res1[9171]);
multi_7x28 multi_7x28_mod_9172(clk,rst,matrix_A[9172],matrix_B[172],mul_res1[9172]);
multi_7x28 multi_7x28_mod_9173(clk,rst,matrix_A[9173],matrix_B[173],mul_res1[9173]);
multi_7x28 multi_7x28_mod_9174(clk,rst,matrix_A[9174],matrix_B[174],mul_res1[9174]);
multi_7x28 multi_7x28_mod_9175(clk,rst,matrix_A[9175],matrix_B[175],mul_res1[9175]);
multi_7x28 multi_7x28_mod_9176(clk,rst,matrix_A[9176],matrix_B[176],mul_res1[9176]);
multi_7x28 multi_7x28_mod_9177(clk,rst,matrix_A[9177],matrix_B[177],mul_res1[9177]);
multi_7x28 multi_7x28_mod_9178(clk,rst,matrix_A[9178],matrix_B[178],mul_res1[9178]);
multi_7x28 multi_7x28_mod_9179(clk,rst,matrix_A[9179],matrix_B[179],mul_res1[9179]);
multi_7x28 multi_7x28_mod_9180(clk,rst,matrix_A[9180],matrix_B[180],mul_res1[9180]);
multi_7x28 multi_7x28_mod_9181(clk,rst,matrix_A[9181],matrix_B[181],mul_res1[9181]);
multi_7x28 multi_7x28_mod_9182(clk,rst,matrix_A[9182],matrix_B[182],mul_res1[9182]);
multi_7x28 multi_7x28_mod_9183(clk,rst,matrix_A[9183],matrix_B[183],mul_res1[9183]);
multi_7x28 multi_7x28_mod_9184(clk,rst,matrix_A[9184],matrix_B[184],mul_res1[9184]);
multi_7x28 multi_7x28_mod_9185(clk,rst,matrix_A[9185],matrix_B[185],mul_res1[9185]);
multi_7x28 multi_7x28_mod_9186(clk,rst,matrix_A[9186],matrix_B[186],mul_res1[9186]);
multi_7x28 multi_7x28_mod_9187(clk,rst,matrix_A[9187],matrix_B[187],mul_res1[9187]);
multi_7x28 multi_7x28_mod_9188(clk,rst,matrix_A[9188],matrix_B[188],mul_res1[9188]);
multi_7x28 multi_7x28_mod_9189(clk,rst,matrix_A[9189],matrix_B[189],mul_res1[9189]);
multi_7x28 multi_7x28_mod_9190(clk,rst,matrix_A[9190],matrix_B[190],mul_res1[9190]);
multi_7x28 multi_7x28_mod_9191(clk,rst,matrix_A[9191],matrix_B[191],mul_res1[9191]);
multi_7x28 multi_7x28_mod_9192(clk,rst,matrix_A[9192],matrix_B[192],mul_res1[9192]);
multi_7x28 multi_7x28_mod_9193(clk,rst,matrix_A[9193],matrix_B[193],mul_res1[9193]);
multi_7x28 multi_7x28_mod_9194(clk,rst,matrix_A[9194],matrix_B[194],mul_res1[9194]);
multi_7x28 multi_7x28_mod_9195(clk,rst,matrix_A[9195],matrix_B[195],mul_res1[9195]);
multi_7x28 multi_7x28_mod_9196(clk,rst,matrix_A[9196],matrix_B[196],mul_res1[9196]);
multi_7x28 multi_7x28_mod_9197(clk,rst,matrix_A[9197],matrix_B[197],mul_res1[9197]);
multi_7x28 multi_7x28_mod_9198(clk,rst,matrix_A[9198],matrix_B[198],mul_res1[9198]);
multi_7x28 multi_7x28_mod_9199(clk,rst,matrix_A[9199],matrix_B[199],mul_res1[9199]);
multi_7x28 multi_7x28_mod_9200(clk,rst,matrix_A[9200],matrix_B[0],mul_res1[9200]);
multi_7x28 multi_7x28_mod_9201(clk,rst,matrix_A[9201],matrix_B[1],mul_res1[9201]);
multi_7x28 multi_7x28_mod_9202(clk,rst,matrix_A[9202],matrix_B[2],mul_res1[9202]);
multi_7x28 multi_7x28_mod_9203(clk,rst,matrix_A[9203],matrix_B[3],mul_res1[9203]);
multi_7x28 multi_7x28_mod_9204(clk,rst,matrix_A[9204],matrix_B[4],mul_res1[9204]);
multi_7x28 multi_7x28_mod_9205(clk,rst,matrix_A[9205],matrix_B[5],mul_res1[9205]);
multi_7x28 multi_7x28_mod_9206(clk,rst,matrix_A[9206],matrix_B[6],mul_res1[9206]);
multi_7x28 multi_7x28_mod_9207(clk,rst,matrix_A[9207],matrix_B[7],mul_res1[9207]);
multi_7x28 multi_7x28_mod_9208(clk,rst,matrix_A[9208],matrix_B[8],mul_res1[9208]);
multi_7x28 multi_7x28_mod_9209(clk,rst,matrix_A[9209],matrix_B[9],mul_res1[9209]);
multi_7x28 multi_7x28_mod_9210(clk,rst,matrix_A[9210],matrix_B[10],mul_res1[9210]);
multi_7x28 multi_7x28_mod_9211(clk,rst,matrix_A[9211],matrix_B[11],mul_res1[9211]);
multi_7x28 multi_7x28_mod_9212(clk,rst,matrix_A[9212],matrix_B[12],mul_res1[9212]);
multi_7x28 multi_7x28_mod_9213(clk,rst,matrix_A[9213],matrix_B[13],mul_res1[9213]);
multi_7x28 multi_7x28_mod_9214(clk,rst,matrix_A[9214],matrix_B[14],mul_res1[9214]);
multi_7x28 multi_7x28_mod_9215(clk,rst,matrix_A[9215],matrix_B[15],mul_res1[9215]);
multi_7x28 multi_7x28_mod_9216(clk,rst,matrix_A[9216],matrix_B[16],mul_res1[9216]);
multi_7x28 multi_7x28_mod_9217(clk,rst,matrix_A[9217],matrix_B[17],mul_res1[9217]);
multi_7x28 multi_7x28_mod_9218(clk,rst,matrix_A[9218],matrix_B[18],mul_res1[9218]);
multi_7x28 multi_7x28_mod_9219(clk,rst,matrix_A[9219],matrix_B[19],mul_res1[9219]);
multi_7x28 multi_7x28_mod_9220(clk,rst,matrix_A[9220],matrix_B[20],mul_res1[9220]);
multi_7x28 multi_7x28_mod_9221(clk,rst,matrix_A[9221],matrix_B[21],mul_res1[9221]);
multi_7x28 multi_7x28_mod_9222(clk,rst,matrix_A[9222],matrix_B[22],mul_res1[9222]);
multi_7x28 multi_7x28_mod_9223(clk,rst,matrix_A[9223],matrix_B[23],mul_res1[9223]);
multi_7x28 multi_7x28_mod_9224(clk,rst,matrix_A[9224],matrix_B[24],mul_res1[9224]);
multi_7x28 multi_7x28_mod_9225(clk,rst,matrix_A[9225],matrix_B[25],mul_res1[9225]);
multi_7x28 multi_7x28_mod_9226(clk,rst,matrix_A[9226],matrix_B[26],mul_res1[9226]);
multi_7x28 multi_7x28_mod_9227(clk,rst,matrix_A[9227],matrix_B[27],mul_res1[9227]);
multi_7x28 multi_7x28_mod_9228(clk,rst,matrix_A[9228],matrix_B[28],mul_res1[9228]);
multi_7x28 multi_7x28_mod_9229(clk,rst,matrix_A[9229],matrix_B[29],mul_res1[9229]);
multi_7x28 multi_7x28_mod_9230(clk,rst,matrix_A[9230],matrix_B[30],mul_res1[9230]);
multi_7x28 multi_7x28_mod_9231(clk,rst,matrix_A[9231],matrix_B[31],mul_res1[9231]);
multi_7x28 multi_7x28_mod_9232(clk,rst,matrix_A[9232],matrix_B[32],mul_res1[9232]);
multi_7x28 multi_7x28_mod_9233(clk,rst,matrix_A[9233],matrix_B[33],mul_res1[9233]);
multi_7x28 multi_7x28_mod_9234(clk,rst,matrix_A[9234],matrix_B[34],mul_res1[9234]);
multi_7x28 multi_7x28_mod_9235(clk,rst,matrix_A[9235],matrix_B[35],mul_res1[9235]);
multi_7x28 multi_7x28_mod_9236(clk,rst,matrix_A[9236],matrix_B[36],mul_res1[9236]);
multi_7x28 multi_7x28_mod_9237(clk,rst,matrix_A[9237],matrix_B[37],mul_res1[9237]);
multi_7x28 multi_7x28_mod_9238(clk,rst,matrix_A[9238],matrix_B[38],mul_res1[9238]);
multi_7x28 multi_7x28_mod_9239(clk,rst,matrix_A[9239],matrix_B[39],mul_res1[9239]);
multi_7x28 multi_7x28_mod_9240(clk,rst,matrix_A[9240],matrix_B[40],mul_res1[9240]);
multi_7x28 multi_7x28_mod_9241(clk,rst,matrix_A[9241],matrix_B[41],mul_res1[9241]);
multi_7x28 multi_7x28_mod_9242(clk,rst,matrix_A[9242],matrix_B[42],mul_res1[9242]);
multi_7x28 multi_7x28_mod_9243(clk,rst,matrix_A[9243],matrix_B[43],mul_res1[9243]);
multi_7x28 multi_7x28_mod_9244(clk,rst,matrix_A[9244],matrix_B[44],mul_res1[9244]);
multi_7x28 multi_7x28_mod_9245(clk,rst,matrix_A[9245],matrix_B[45],mul_res1[9245]);
multi_7x28 multi_7x28_mod_9246(clk,rst,matrix_A[9246],matrix_B[46],mul_res1[9246]);
multi_7x28 multi_7x28_mod_9247(clk,rst,matrix_A[9247],matrix_B[47],mul_res1[9247]);
multi_7x28 multi_7x28_mod_9248(clk,rst,matrix_A[9248],matrix_B[48],mul_res1[9248]);
multi_7x28 multi_7x28_mod_9249(clk,rst,matrix_A[9249],matrix_B[49],mul_res1[9249]);
multi_7x28 multi_7x28_mod_9250(clk,rst,matrix_A[9250],matrix_B[50],mul_res1[9250]);
multi_7x28 multi_7x28_mod_9251(clk,rst,matrix_A[9251],matrix_B[51],mul_res1[9251]);
multi_7x28 multi_7x28_mod_9252(clk,rst,matrix_A[9252],matrix_B[52],mul_res1[9252]);
multi_7x28 multi_7x28_mod_9253(clk,rst,matrix_A[9253],matrix_B[53],mul_res1[9253]);
multi_7x28 multi_7x28_mod_9254(clk,rst,matrix_A[9254],matrix_B[54],mul_res1[9254]);
multi_7x28 multi_7x28_mod_9255(clk,rst,matrix_A[9255],matrix_B[55],mul_res1[9255]);
multi_7x28 multi_7x28_mod_9256(clk,rst,matrix_A[9256],matrix_B[56],mul_res1[9256]);
multi_7x28 multi_7x28_mod_9257(clk,rst,matrix_A[9257],matrix_B[57],mul_res1[9257]);
multi_7x28 multi_7x28_mod_9258(clk,rst,matrix_A[9258],matrix_B[58],mul_res1[9258]);
multi_7x28 multi_7x28_mod_9259(clk,rst,matrix_A[9259],matrix_B[59],mul_res1[9259]);
multi_7x28 multi_7x28_mod_9260(clk,rst,matrix_A[9260],matrix_B[60],mul_res1[9260]);
multi_7x28 multi_7x28_mod_9261(clk,rst,matrix_A[9261],matrix_B[61],mul_res1[9261]);
multi_7x28 multi_7x28_mod_9262(clk,rst,matrix_A[9262],matrix_B[62],mul_res1[9262]);
multi_7x28 multi_7x28_mod_9263(clk,rst,matrix_A[9263],matrix_B[63],mul_res1[9263]);
multi_7x28 multi_7x28_mod_9264(clk,rst,matrix_A[9264],matrix_B[64],mul_res1[9264]);
multi_7x28 multi_7x28_mod_9265(clk,rst,matrix_A[9265],matrix_B[65],mul_res1[9265]);
multi_7x28 multi_7x28_mod_9266(clk,rst,matrix_A[9266],matrix_B[66],mul_res1[9266]);
multi_7x28 multi_7x28_mod_9267(clk,rst,matrix_A[9267],matrix_B[67],mul_res1[9267]);
multi_7x28 multi_7x28_mod_9268(clk,rst,matrix_A[9268],matrix_B[68],mul_res1[9268]);
multi_7x28 multi_7x28_mod_9269(clk,rst,matrix_A[9269],matrix_B[69],mul_res1[9269]);
multi_7x28 multi_7x28_mod_9270(clk,rst,matrix_A[9270],matrix_B[70],mul_res1[9270]);
multi_7x28 multi_7x28_mod_9271(clk,rst,matrix_A[9271],matrix_B[71],mul_res1[9271]);
multi_7x28 multi_7x28_mod_9272(clk,rst,matrix_A[9272],matrix_B[72],mul_res1[9272]);
multi_7x28 multi_7x28_mod_9273(clk,rst,matrix_A[9273],matrix_B[73],mul_res1[9273]);
multi_7x28 multi_7x28_mod_9274(clk,rst,matrix_A[9274],matrix_B[74],mul_res1[9274]);
multi_7x28 multi_7x28_mod_9275(clk,rst,matrix_A[9275],matrix_B[75],mul_res1[9275]);
multi_7x28 multi_7x28_mod_9276(clk,rst,matrix_A[9276],matrix_B[76],mul_res1[9276]);
multi_7x28 multi_7x28_mod_9277(clk,rst,matrix_A[9277],matrix_B[77],mul_res1[9277]);
multi_7x28 multi_7x28_mod_9278(clk,rst,matrix_A[9278],matrix_B[78],mul_res1[9278]);
multi_7x28 multi_7x28_mod_9279(clk,rst,matrix_A[9279],matrix_B[79],mul_res1[9279]);
multi_7x28 multi_7x28_mod_9280(clk,rst,matrix_A[9280],matrix_B[80],mul_res1[9280]);
multi_7x28 multi_7x28_mod_9281(clk,rst,matrix_A[9281],matrix_B[81],mul_res1[9281]);
multi_7x28 multi_7x28_mod_9282(clk,rst,matrix_A[9282],matrix_B[82],mul_res1[9282]);
multi_7x28 multi_7x28_mod_9283(clk,rst,matrix_A[9283],matrix_B[83],mul_res1[9283]);
multi_7x28 multi_7x28_mod_9284(clk,rst,matrix_A[9284],matrix_B[84],mul_res1[9284]);
multi_7x28 multi_7x28_mod_9285(clk,rst,matrix_A[9285],matrix_B[85],mul_res1[9285]);
multi_7x28 multi_7x28_mod_9286(clk,rst,matrix_A[9286],matrix_B[86],mul_res1[9286]);
multi_7x28 multi_7x28_mod_9287(clk,rst,matrix_A[9287],matrix_B[87],mul_res1[9287]);
multi_7x28 multi_7x28_mod_9288(clk,rst,matrix_A[9288],matrix_B[88],mul_res1[9288]);
multi_7x28 multi_7x28_mod_9289(clk,rst,matrix_A[9289],matrix_B[89],mul_res1[9289]);
multi_7x28 multi_7x28_mod_9290(clk,rst,matrix_A[9290],matrix_B[90],mul_res1[9290]);
multi_7x28 multi_7x28_mod_9291(clk,rst,matrix_A[9291],matrix_B[91],mul_res1[9291]);
multi_7x28 multi_7x28_mod_9292(clk,rst,matrix_A[9292],matrix_B[92],mul_res1[9292]);
multi_7x28 multi_7x28_mod_9293(clk,rst,matrix_A[9293],matrix_B[93],mul_res1[9293]);
multi_7x28 multi_7x28_mod_9294(clk,rst,matrix_A[9294],matrix_B[94],mul_res1[9294]);
multi_7x28 multi_7x28_mod_9295(clk,rst,matrix_A[9295],matrix_B[95],mul_res1[9295]);
multi_7x28 multi_7x28_mod_9296(clk,rst,matrix_A[9296],matrix_B[96],mul_res1[9296]);
multi_7x28 multi_7x28_mod_9297(clk,rst,matrix_A[9297],matrix_B[97],mul_res1[9297]);
multi_7x28 multi_7x28_mod_9298(clk,rst,matrix_A[9298],matrix_B[98],mul_res1[9298]);
multi_7x28 multi_7x28_mod_9299(clk,rst,matrix_A[9299],matrix_B[99],mul_res1[9299]);
multi_7x28 multi_7x28_mod_9300(clk,rst,matrix_A[9300],matrix_B[100],mul_res1[9300]);
multi_7x28 multi_7x28_mod_9301(clk,rst,matrix_A[9301],matrix_B[101],mul_res1[9301]);
multi_7x28 multi_7x28_mod_9302(clk,rst,matrix_A[9302],matrix_B[102],mul_res1[9302]);
multi_7x28 multi_7x28_mod_9303(clk,rst,matrix_A[9303],matrix_B[103],mul_res1[9303]);
multi_7x28 multi_7x28_mod_9304(clk,rst,matrix_A[9304],matrix_B[104],mul_res1[9304]);
multi_7x28 multi_7x28_mod_9305(clk,rst,matrix_A[9305],matrix_B[105],mul_res1[9305]);
multi_7x28 multi_7x28_mod_9306(clk,rst,matrix_A[9306],matrix_B[106],mul_res1[9306]);
multi_7x28 multi_7x28_mod_9307(clk,rst,matrix_A[9307],matrix_B[107],mul_res1[9307]);
multi_7x28 multi_7x28_mod_9308(clk,rst,matrix_A[9308],matrix_B[108],mul_res1[9308]);
multi_7x28 multi_7x28_mod_9309(clk,rst,matrix_A[9309],matrix_B[109],mul_res1[9309]);
multi_7x28 multi_7x28_mod_9310(clk,rst,matrix_A[9310],matrix_B[110],mul_res1[9310]);
multi_7x28 multi_7x28_mod_9311(clk,rst,matrix_A[9311],matrix_B[111],mul_res1[9311]);
multi_7x28 multi_7x28_mod_9312(clk,rst,matrix_A[9312],matrix_B[112],mul_res1[9312]);
multi_7x28 multi_7x28_mod_9313(clk,rst,matrix_A[9313],matrix_B[113],mul_res1[9313]);
multi_7x28 multi_7x28_mod_9314(clk,rst,matrix_A[9314],matrix_B[114],mul_res1[9314]);
multi_7x28 multi_7x28_mod_9315(clk,rst,matrix_A[9315],matrix_B[115],mul_res1[9315]);
multi_7x28 multi_7x28_mod_9316(clk,rst,matrix_A[9316],matrix_B[116],mul_res1[9316]);
multi_7x28 multi_7x28_mod_9317(clk,rst,matrix_A[9317],matrix_B[117],mul_res1[9317]);
multi_7x28 multi_7x28_mod_9318(clk,rst,matrix_A[9318],matrix_B[118],mul_res1[9318]);
multi_7x28 multi_7x28_mod_9319(clk,rst,matrix_A[9319],matrix_B[119],mul_res1[9319]);
multi_7x28 multi_7x28_mod_9320(clk,rst,matrix_A[9320],matrix_B[120],mul_res1[9320]);
multi_7x28 multi_7x28_mod_9321(clk,rst,matrix_A[9321],matrix_B[121],mul_res1[9321]);
multi_7x28 multi_7x28_mod_9322(clk,rst,matrix_A[9322],matrix_B[122],mul_res1[9322]);
multi_7x28 multi_7x28_mod_9323(clk,rst,matrix_A[9323],matrix_B[123],mul_res1[9323]);
multi_7x28 multi_7x28_mod_9324(clk,rst,matrix_A[9324],matrix_B[124],mul_res1[9324]);
multi_7x28 multi_7x28_mod_9325(clk,rst,matrix_A[9325],matrix_B[125],mul_res1[9325]);
multi_7x28 multi_7x28_mod_9326(clk,rst,matrix_A[9326],matrix_B[126],mul_res1[9326]);
multi_7x28 multi_7x28_mod_9327(clk,rst,matrix_A[9327],matrix_B[127],mul_res1[9327]);
multi_7x28 multi_7x28_mod_9328(clk,rst,matrix_A[9328],matrix_B[128],mul_res1[9328]);
multi_7x28 multi_7x28_mod_9329(clk,rst,matrix_A[9329],matrix_B[129],mul_res1[9329]);
multi_7x28 multi_7x28_mod_9330(clk,rst,matrix_A[9330],matrix_B[130],mul_res1[9330]);
multi_7x28 multi_7x28_mod_9331(clk,rst,matrix_A[9331],matrix_B[131],mul_res1[9331]);
multi_7x28 multi_7x28_mod_9332(clk,rst,matrix_A[9332],matrix_B[132],mul_res1[9332]);
multi_7x28 multi_7x28_mod_9333(clk,rst,matrix_A[9333],matrix_B[133],mul_res1[9333]);
multi_7x28 multi_7x28_mod_9334(clk,rst,matrix_A[9334],matrix_B[134],mul_res1[9334]);
multi_7x28 multi_7x28_mod_9335(clk,rst,matrix_A[9335],matrix_B[135],mul_res1[9335]);
multi_7x28 multi_7x28_mod_9336(clk,rst,matrix_A[9336],matrix_B[136],mul_res1[9336]);
multi_7x28 multi_7x28_mod_9337(clk,rst,matrix_A[9337],matrix_B[137],mul_res1[9337]);
multi_7x28 multi_7x28_mod_9338(clk,rst,matrix_A[9338],matrix_B[138],mul_res1[9338]);
multi_7x28 multi_7x28_mod_9339(clk,rst,matrix_A[9339],matrix_B[139],mul_res1[9339]);
multi_7x28 multi_7x28_mod_9340(clk,rst,matrix_A[9340],matrix_B[140],mul_res1[9340]);
multi_7x28 multi_7x28_mod_9341(clk,rst,matrix_A[9341],matrix_B[141],mul_res1[9341]);
multi_7x28 multi_7x28_mod_9342(clk,rst,matrix_A[9342],matrix_B[142],mul_res1[9342]);
multi_7x28 multi_7x28_mod_9343(clk,rst,matrix_A[9343],matrix_B[143],mul_res1[9343]);
multi_7x28 multi_7x28_mod_9344(clk,rst,matrix_A[9344],matrix_B[144],mul_res1[9344]);
multi_7x28 multi_7x28_mod_9345(clk,rst,matrix_A[9345],matrix_B[145],mul_res1[9345]);
multi_7x28 multi_7x28_mod_9346(clk,rst,matrix_A[9346],matrix_B[146],mul_res1[9346]);
multi_7x28 multi_7x28_mod_9347(clk,rst,matrix_A[9347],matrix_B[147],mul_res1[9347]);
multi_7x28 multi_7x28_mod_9348(clk,rst,matrix_A[9348],matrix_B[148],mul_res1[9348]);
multi_7x28 multi_7x28_mod_9349(clk,rst,matrix_A[9349],matrix_B[149],mul_res1[9349]);
multi_7x28 multi_7x28_mod_9350(clk,rst,matrix_A[9350],matrix_B[150],mul_res1[9350]);
multi_7x28 multi_7x28_mod_9351(clk,rst,matrix_A[9351],matrix_B[151],mul_res1[9351]);
multi_7x28 multi_7x28_mod_9352(clk,rst,matrix_A[9352],matrix_B[152],mul_res1[9352]);
multi_7x28 multi_7x28_mod_9353(clk,rst,matrix_A[9353],matrix_B[153],mul_res1[9353]);
multi_7x28 multi_7x28_mod_9354(clk,rst,matrix_A[9354],matrix_B[154],mul_res1[9354]);
multi_7x28 multi_7x28_mod_9355(clk,rst,matrix_A[9355],matrix_B[155],mul_res1[9355]);
multi_7x28 multi_7x28_mod_9356(clk,rst,matrix_A[9356],matrix_B[156],mul_res1[9356]);
multi_7x28 multi_7x28_mod_9357(clk,rst,matrix_A[9357],matrix_B[157],mul_res1[9357]);
multi_7x28 multi_7x28_mod_9358(clk,rst,matrix_A[9358],matrix_B[158],mul_res1[9358]);
multi_7x28 multi_7x28_mod_9359(clk,rst,matrix_A[9359],matrix_B[159],mul_res1[9359]);
multi_7x28 multi_7x28_mod_9360(clk,rst,matrix_A[9360],matrix_B[160],mul_res1[9360]);
multi_7x28 multi_7x28_mod_9361(clk,rst,matrix_A[9361],matrix_B[161],mul_res1[9361]);
multi_7x28 multi_7x28_mod_9362(clk,rst,matrix_A[9362],matrix_B[162],mul_res1[9362]);
multi_7x28 multi_7x28_mod_9363(clk,rst,matrix_A[9363],matrix_B[163],mul_res1[9363]);
multi_7x28 multi_7x28_mod_9364(clk,rst,matrix_A[9364],matrix_B[164],mul_res1[9364]);
multi_7x28 multi_7x28_mod_9365(clk,rst,matrix_A[9365],matrix_B[165],mul_res1[9365]);
multi_7x28 multi_7x28_mod_9366(clk,rst,matrix_A[9366],matrix_B[166],mul_res1[9366]);
multi_7x28 multi_7x28_mod_9367(clk,rst,matrix_A[9367],matrix_B[167],mul_res1[9367]);
multi_7x28 multi_7x28_mod_9368(clk,rst,matrix_A[9368],matrix_B[168],mul_res1[9368]);
multi_7x28 multi_7x28_mod_9369(clk,rst,matrix_A[9369],matrix_B[169],mul_res1[9369]);
multi_7x28 multi_7x28_mod_9370(clk,rst,matrix_A[9370],matrix_B[170],mul_res1[9370]);
multi_7x28 multi_7x28_mod_9371(clk,rst,matrix_A[9371],matrix_B[171],mul_res1[9371]);
multi_7x28 multi_7x28_mod_9372(clk,rst,matrix_A[9372],matrix_B[172],mul_res1[9372]);
multi_7x28 multi_7x28_mod_9373(clk,rst,matrix_A[9373],matrix_B[173],mul_res1[9373]);
multi_7x28 multi_7x28_mod_9374(clk,rst,matrix_A[9374],matrix_B[174],mul_res1[9374]);
multi_7x28 multi_7x28_mod_9375(clk,rst,matrix_A[9375],matrix_B[175],mul_res1[9375]);
multi_7x28 multi_7x28_mod_9376(clk,rst,matrix_A[9376],matrix_B[176],mul_res1[9376]);
multi_7x28 multi_7x28_mod_9377(clk,rst,matrix_A[9377],matrix_B[177],mul_res1[9377]);
multi_7x28 multi_7x28_mod_9378(clk,rst,matrix_A[9378],matrix_B[178],mul_res1[9378]);
multi_7x28 multi_7x28_mod_9379(clk,rst,matrix_A[9379],matrix_B[179],mul_res1[9379]);
multi_7x28 multi_7x28_mod_9380(clk,rst,matrix_A[9380],matrix_B[180],mul_res1[9380]);
multi_7x28 multi_7x28_mod_9381(clk,rst,matrix_A[9381],matrix_B[181],mul_res1[9381]);
multi_7x28 multi_7x28_mod_9382(clk,rst,matrix_A[9382],matrix_B[182],mul_res1[9382]);
multi_7x28 multi_7x28_mod_9383(clk,rst,matrix_A[9383],matrix_B[183],mul_res1[9383]);
multi_7x28 multi_7x28_mod_9384(clk,rst,matrix_A[9384],matrix_B[184],mul_res1[9384]);
multi_7x28 multi_7x28_mod_9385(clk,rst,matrix_A[9385],matrix_B[185],mul_res1[9385]);
multi_7x28 multi_7x28_mod_9386(clk,rst,matrix_A[9386],matrix_B[186],mul_res1[9386]);
multi_7x28 multi_7x28_mod_9387(clk,rst,matrix_A[9387],matrix_B[187],mul_res1[9387]);
multi_7x28 multi_7x28_mod_9388(clk,rst,matrix_A[9388],matrix_B[188],mul_res1[9388]);
multi_7x28 multi_7x28_mod_9389(clk,rst,matrix_A[9389],matrix_B[189],mul_res1[9389]);
multi_7x28 multi_7x28_mod_9390(clk,rst,matrix_A[9390],matrix_B[190],mul_res1[9390]);
multi_7x28 multi_7x28_mod_9391(clk,rst,matrix_A[9391],matrix_B[191],mul_res1[9391]);
multi_7x28 multi_7x28_mod_9392(clk,rst,matrix_A[9392],matrix_B[192],mul_res1[9392]);
multi_7x28 multi_7x28_mod_9393(clk,rst,matrix_A[9393],matrix_B[193],mul_res1[9393]);
multi_7x28 multi_7x28_mod_9394(clk,rst,matrix_A[9394],matrix_B[194],mul_res1[9394]);
multi_7x28 multi_7x28_mod_9395(clk,rst,matrix_A[9395],matrix_B[195],mul_res1[9395]);
multi_7x28 multi_7x28_mod_9396(clk,rst,matrix_A[9396],matrix_B[196],mul_res1[9396]);
multi_7x28 multi_7x28_mod_9397(clk,rst,matrix_A[9397],matrix_B[197],mul_res1[9397]);
multi_7x28 multi_7x28_mod_9398(clk,rst,matrix_A[9398],matrix_B[198],mul_res1[9398]);
multi_7x28 multi_7x28_mod_9399(clk,rst,matrix_A[9399],matrix_B[199],mul_res1[9399]);
multi_7x28 multi_7x28_mod_9400(clk,rst,matrix_A[9400],matrix_B[0],mul_res1[9400]);
multi_7x28 multi_7x28_mod_9401(clk,rst,matrix_A[9401],matrix_B[1],mul_res1[9401]);
multi_7x28 multi_7x28_mod_9402(clk,rst,matrix_A[9402],matrix_B[2],mul_res1[9402]);
multi_7x28 multi_7x28_mod_9403(clk,rst,matrix_A[9403],matrix_B[3],mul_res1[9403]);
multi_7x28 multi_7x28_mod_9404(clk,rst,matrix_A[9404],matrix_B[4],mul_res1[9404]);
multi_7x28 multi_7x28_mod_9405(clk,rst,matrix_A[9405],matrix_B[5],mul_res1[9405]);
multi_7x28 multi_7x28_mod_9406(clk,rst,matrix_A[9406],matrix_B[6],mul_res1[9406]);
multi_7x28 multi_7x28_mod_9407(clk,rst,matrix_A[9407],matrix_B[7],mul_res1[9407]);
multi_7x28 multi_7x28_mod_9408(clk,rst,matrix_A[9408],matrix_B[8],mul_res1[9408]);
multi_7x28 multi_7x28_mod_9409(clk,rst,matrix_A[9409],matrix_B[9],mul_res1[9409]);
multi_7x28 multi_7x28_mod_9410(clk,rst,matrix_A[9410],matrix_B[10],mul_res1[9410]);
multi_7x28 multi_7x28_mod_9411(clk,rst,matrix_A[9411],matrix_B[11],mul_res1[9411]);
multi_7x28 multi_7x28_mod_9412(clk,rst,matrix_A[9412],matrix_B[12],mul_res1[9412]);
multi_7x28 multi_7x28_mod_9413(clk,rst,matrix_A[9413],matrix_B[13],mul_res1[9413]);
multi_7x28 multi_7x28_mod_9414(clk,rst,matrix_A[9414],matrix_B[14],mul_res1[9414]);
multi_7x28 multi_7x28_mod_9415(clk,rst,matrix_A[9415],matrix_B[15],mul_res1[9415]);
multi_7x28 multi_7x28_mod_9416(clk,rst,matrix_A[9416],matrix_B[16],mul_res1[9416]);
multi_7x28 multi_7x28_mod_9417(clk,rst,matrix_A[9417],matrix_B[17],mul_res1[9417]);
multi_7x28 multi_7x28_mod_9418(clk,rst,matrix_A[9418],matrix_B[18],mul_res1[9418]);
multi_7x28 multi_7x28_mod_9419(clk,rst,matrix_A[9419],matrix_B[19],mul_res1[9419]);
multi_7x28 multi_7x28_mod_9420(clk,rst,matrix_A[9420],matrix_B[20],mul_res1[9420]);
multi_7x28 multi_7x28_mod_9421(clk,rst,matrix_A[9421],matrix_B[21],mul_res1[9421]);
multi_7x28 multi_7x28_mod_9422(clk,rst,matrix_A[9422],matrix_B[22],mul_res1[9422]);
multi_7x28 multi_7x28_mod_9423(clk,rst,matrix_A[9423],matrix_B[23],mul_res1[9423]);
multi_7x28 multi_7x28_mod_9424(clk,rst,matrix_A[9424],matrix_B[24],mul_res1[9424]);
multi_7x28 multi_7x28_mod_9425(clk,rst,matrix_A[9425],matrix_B[25],mul_res1[9425]);
multi_7x28 multi_7x28_mod_9426(clk,rst,matrix_A[9426],matrix_B[26],mul_res1[9426]);
multi_7x28 multi_7x28_mod_9427(clk,rst,matrix_A[9427],matrix_B[27],mul_res1[9427]);
multi_7x28 multi_7x28_mod_9428(clk,rst,matrix_A[9428],matrix_B[28],mul_res1[9428]);
multi_7x28 multi_7x28_mod_9429(clk,rst,matrix_A[9429],matrix_B[29],mul_res1[9429]);
multi_7x28 multi_7x28_mod_9430(clk,rst,matrix_A[9430],matrix_B[30],mul_res1[9430]);
multi_7x28 multi_7x28_mod_9431(clk,rst,matrix_A[9431],matrix_B[31],mul_res1[9431]);
multi_7x28 multi_7x28_mod_9432(clk,rst,matrix_A[9432],matrix_B[32],mul_res1[9432]);
multi_7x28 multi_7x28_mod_9433(clk,rst,matrix_A[9433],matrix_B[33],mul_res1[9433]);
multi_7x28 multi_7x28_mod_9434(clk,rst,matrix_A[9434],matrix_B[34],mul_res1[9434]);
multi_7x28 multi_7x28_mod_9435(clk,rst,matrix_A[9435],matrix_B[35],mul_res1[9435]);
multi_7x28 multi_7x28_mod_9436(clk,rst,matrix_A[9436],matrix_B[36],mul_res1[9436]);
multi_7x28 multi_7x28_mod_9437(clk,rst,matrix_A[9437],matrix_B[37],mul_res1[9437]);
multi_7x28 multi_7x28_mod_9438(clk,rst,matrix_A[9438],matrix_B[38],mul_res1[9438]);
multi_7x28 multi_7x28_mod_9439(clk,rst,matrix_A[9439],matrix_B[39],mul_res1[9439]);
multi_7x28 multi_7x28_mod_9440(clk,rst,matrix_A[9440],matrix_B[40],mul_res1[9440]);
multi_7x28 multi_7x28_mod_9441(clk,rst,matrix_A[9441],matrix_B[41],mul_res1[9441]);
multi_7x28 multi_7x28_mod_9442(clk,rst,matrix_A[9442],matrix_B[42],mul_res1[9442]);
multi_7x28 multi_7x28_mod_9443(clk,rst,matrix_A[9443],matrix_B[43],mul_res1[9443]);
multi_7x28 multi_7x28_mod_9444(clk,rst,matrix_A[9444],matrix_B[44],mul_res1[9444]);
multi_7x28 multi_7x28_mod_9445(clk,rst,matrix_A[9445],matrix_B[45],mul_res1[9445]);
multi_7x28 multi_7x28_mod_9446(clk,rst,matrix_A[9446],matrix_B[46],mul_res1[9446]);
multi_7x28 multi_7x28_mod_9447(clk,rst,matrix_A[9447],matrix_B[47],mul_res1[9447]);
multi_7x28 multi_7x28_mod_9448(clk,rst,matrix_A[9448],matrix_B[48],mul_res1[9448]);
multi_7x28 multi_7x28_mod_9449(clk,rst,matrix_A[9449],matrix_B[49],mul_res1[9449]);
multi_7x28 multi_7x28_mod_9450(clk,rst,matrix_A[9450],matrix_B[50],mul_res1[9450]);
multi_7x28 multi_7x28_mod_9451(clk,rst,matrix_A[9451],matrix_B[51],mul_res1[9451]);
multi_7x28 multi_7x28_mod_9452(clk,rst,matrix_A[9452],matrix_B[52],mul_res1[9452]);
multi_7x28 multi_7x28_mod_9453(clk,rst,matrix_A[9453],matrix_B[53],mul_res1[9453]);
multi_7x28 multi_7x28_mod_9454(clk,rst,matrix_A[9454],matrix_B[54],mul_res1[9454]);
multi_7x28 multi_7x28_mod_9455(clk,rst,matrix_A[9455],matrix_B[55],mul_res1[9455]);
multi_7x28 multi_7x28_mod_9456(clk,rst,matrix_A[9456],matrix_B[56],mul_res1[9456]);
multi_7x28 multi_7x28_mod_9457(clk,rst,matrix_A[9457],matrix_B[57],mul_res1[9457]);
multi_7x28 multi_7x28_mod_9458(clk,rst,matrix_A[9458],matrix_B[58],mul_res1[9458]);
multi_7x28 multi_7x28_mod_9459(clk,rst,matrix_A[9459],matrix_B[59],mul_res1[9459]);
multi_7x28 multi_7x28_mod_9460(clk,rst,matrix_A[9460],matrix_B[60],mul_res1[9460]);
multi_7x28 multi_7x28_mod_9461(clk,rst,matrix_A[9461],matrix_B[61],mul_res1[9461]);
multi_7x28 multi_7x28_mod_9462(clk,rst,matrix_A[9462],matrix_B[62],mul_res1[9462]);
multi_7x28 multi_7x28_mod_9463(clk,rst,matrix_A[9463],matrix_B[63],mul_res1[9463]);
multi_7x28 multi_7x28_mod_9464(clk,rst,matrix_A[9464],matrix_B[64],mul_res1[9464]);
multi_7x28 multi_7x28_mod_9465(clk,rst,matrix_A[9465],matrix_B[65],mul_res1[9465]);
multi_7x28 multi_7x28_mod_9466(clk,rst,matrix_A[9466],matrix_B[66],mul_res1[9466]);
multi_7x28 multi_7x28_mod_9467(clk,rst,matrix_A[9467],matrix_B[67],mul_res1[9467]);
multi_7x28 multi_7x28_mod_9468(clk,rst,matrix_A[9468],matrix_B[68],mul_res1[9468]);
multi_7x28 multi_7x28_mod_9469(clk,rst,matrix_A[9469],matrix_B[69],mul_res1[9469]);
multi_7x28 multi_7x28_mod_9470(clk,rst,matrix_A[9470],matrix_B[70],mul_res1[9470]);
multi_7x28 multi_7x28_mod_9471(clk,rst,matrix_A[9471],matrix_B[71],mul_res1[9471]);
multi_7x28 multi_7x28_mod_9472(clk,rst,matrix_A[9472],matrix_B[72],mul_res1[9472]);
multi_7x28 multi_7x28_mod_9473(clk,rst,matrix_A[9473],matrix_B[73],mul_res1[9473]);
multi_7x28 multi_7x28_mod_9474(clk,rst,matrix_A[9474],matrix_B[74],mul_res1[9474]);
multi_7x28 multi_7x28_mod_9475(clk,rst,matrix_A[9475],matrix_B[75],mul_res1[9475]);
multi_7x28 multi_7x28_mod_9476(clk,rst,matrix_A[9476],matrix_B[76],mul_res1[9476]);
multi_7x28 multi_7x28_mod_9477(clk,rst,matrix_A[9477],matrix_B[77],mul_res1[9477]);
multi_7x28 multi_7x28_mod_9478(clk,rst,matrix_A[9478],matrix_B[78],mul_res1[9478]);
multi_7x28 multi_7x28_mod_9479(clk,rst,matrix_A[9479],matrix_B[79],mul_res1[9479]);
multi_7x28 multi_7x28_mod_9480(clk,rst,matrix_A[9480],matrix_B[80],mul_res1[9480]);
multi_7x28 multi_7x28_mod_9481(clk,rst,matrix_A[9481],matrix_B[81],mul_res1[9481]);
multi_7x28 multi_7x28_mod_9482(clk,rst,matrix_A[9482],matrix_B[82],mul_res1[9482]);
multi_7x28 multi_7x28_mod_9483(clk,rst,matrix_A[9483],matrix_B[83],mul_res1[9483]);
multi_7x28 multi_7x28_mod_9484(clk,rst,matrix_A[9484],matrix_B[84],mul_res1[9484]);
multi_7x28 multi_7x28_mod_9485(clk,rst,matrix_A[9485],matrix_B[85],mul_res1[9485]);
multi_7x28 multi_7x28_mod_9486(clk,rst,matrix_A[9486],matrix_B[86],mul_res1[9486]);
multi_7x28 multi_7x28_mod_9487(clk,rst,matrix_A[9487],matrix_B[87],mul_res1[9487]);
multi_7x28 multi_7x28_mod_9488(clk,rst,matrix_A[9488],matrix_B[88],mul_res1[9488]);
multi_7x28 multi_7x28_mod_9489(clk,rst,matrix_A[9489],matrix_B[89],mul_res1[9489]);
multi_7x28 multi_7x28_mod_9490(clk,rst,matrix_A[9490],matrix_B[90],mul_res1[9490]);
multi_7x28 multi_7x28_mod_9491(clk,rst,matrix_A[9491],matrix_B[91],mul_res1[9491]);
multi_7x28 multi_7x28_mod_9492(clk,rst,matrix_A[9492],matrix_B[92],mul_res1[9492]);
multi_7x28 multi_7x28_mod_9493(clk,rst,matrix_A[9493],matrix_B[93],mul_res1[9493]);
multi_7x28 multi_7x28_mod_9494(clk,rst,matrix_A[9494],matrix_B[94],mul_res1[9494]);
multi_7x28 multi_7x28_mod_9495(clk,rst,matrix_A[9495],matrix_B[95],mul_res1[9495]);
multi_7x28 multi_7x28_mod_9496(clk,rst,matrix_A[9496],matrix_B[96],mul_res1[9496]);
multi_7x28 multi_7x28_mod_9497(clk,rst,matrix_A[9497],matrix_B[97],mul_res1[9497]);
multi_7x28 multi_7x28_mod_9498(clk,rst,matrix_A[9498],matrix_B[98],mul_res1[9498]);
multi_7x28 multi_7x28_mod_9499(clk,rst,matrix_A[9499],matrix_B[99],mul_res1[9499]);
multi_7x28 multi_7x28_mod_9500(clk,rst,matrix_A[9500],matrix_B[100],mul_res1[9500]);
multi_7x28 multi_7x28_mod_9501(clk,rst,matrix_A[9501],matrix_B[101],mul_res1[9501]);
multi_7x28 multi_7x28_mod_9502(clk,rst,matrix_A[9502],matrix_B[102],mul_res1[9502]);
multi_7x28 multi_7x28_mod_9503(clk,rst,matrix_A[9503],matrix_B[103],mul_res1[9503]);
multi_7x28 multi_7x28_mod_9504(clk,rst,matrix_A[9504],matrix_B[104],mul_res1[9504]);
multi_7x28 multi_7x28_mod_9505(clk,rst,matrix_A[9505],matrix_B[105],mul_res1[9505]);
multi_7x28 multi_7x28_mod_9506(clk,rst,matrix_A[9506],matrix_B[106],mul_res1[9506]);
multi_7x28 multi_7x28_mod_9507(clk,rst,matrix_A[9507],matrix_B[107],mul_res1[9507]);
multi_7x28 multi_7x28_mod_9508(clk,rst,matrix_A[9508],matrix_B[108],mul_res1[9508]);
multi_7x28 multi_7x28_mod_9509(clk,rst,matrix_A[9509],matrix_B[109],mul_res1[9509]);
multi_7x28 multi_7x28_mod_9510(clk,rst,matrix_A[9510],matrix_B[110],mul_res1[9510]);
multi_7x28 multi_7x28_mod_9511(clk,rst,matrix_A[9511],matrix_B[111],mul_res1[9511]);
multi_7x28 multi_7x28_mod_9512(clk,rst,matrix_A[9512],matrix_B[112],mul_res1[9512]);
multi_7x28 multi_7x28_mod_9513(clk,rst,matrix_A[9513],matrix_B[113],mul_res1[9513]);
multi_7x28 multi_7x28_mod_9514(clk,rst,matrix_A[9514],matrix_B[114],mul_res1[9514]);
multi_7x28 multi_7x28_mod_9515(clk,rst,matrix_A[9515],matrix_B[115],mul_res1[9515]);
multi_7x28 multi_7x28_mod_9516(clk,rst,matrix_A[9516],matrix_B[116],mul_res1[9516]);
multi_7x28 multi_7x28_mod_9517(clk,rst,matrix_A[9517],matrix_B[117],mul_res1[9517]);
multi_7x28 multi_7x28_mod_9518(clk,rst,matrix_A[9518],matrix_B[118],mul_res1[9518]);
multi_7x28 multi_7x28_mod_9519(clk,rst,matrix_A[9519],matrix_B[119],mul_res1[9519]);
multi_7x28 multi_7x28_mod_9520(clk,rst,matrix_A[9520],matrix_B[120],mul_res1[9520]);
multi_7x28 multi_7x28_mod_9521(clk,rst,matrix_A[9521],matrix_B[121],mul_res1[9521]);
multi_7x28 multi_7x28_mod_9522(clk,rst,matrix_A[9522],matrix_B[122],mul_res1[9522]);
multi_7x28 multi_7x28_mod_9523(clk,rst,matrix_A[9523],matrix_B[123],mul_res1[9523]);
multi_7x28 multi_7x28_mod_9524(clk,rst,matrix_A[9524],matrix_B[124],mul_res1[9524]);
multi_7x28 multi_7x28_mod_9525(clk,rst,matrix_A[9525],matrix_B[125],mul_res1[9525]);
multi_7x28 multi_7x28_mod_9526(clk,rst,matrix_A[9526],matrix_B[126],mul_res1[9526]);
multi_7x28 multi_7x28_mod_9527(clk,rst,matrix_A[9527],matrix_B[127],mul_res1[9527]);
multi_7x28 multi_7x28_mod_9528(clk,rst,matrix_A[9528],matrix_B[128],mul_res1[9528]);
multi_7x28 multi_7x28_mod_9529(clk,rst,matrix_A[9529],matrix_B[129],mul_res1[9529]);
multi_7x28 multi_7x28_mod_9530(clk,rst,matrix_A[9530],matrix_B[130],mul_res1[9530]);
multi_7x28 multi_7x28_mod_9531(clk,rst,matrix_A[9531],matrix_B[131],mul_res1[9531]);
multi_7x28 multi_7x28_mod_9532(clk,rst,matrix_A[9532],matrix_B[132],mul_res1[9532]);
multi_7x28 multi_7x28_mod_9533(clk,rst,matrix_A[9533],matrix_B[133],mul_res1[9533]);
multi_7x28 multi_7x28_mod_9534(clk,rst,matrix_A[9534],matrix_B[134],mul_res1[9534]);
multi_7x28 multi_7x28_mod_9535(clk,rst,matrix_A[9535],matrix_B[135],mul_res1[9535]);
multi_7x28 multi_7x28_mod_9536(clk,rst,matrix_A[9536],matrix_B[136],mul_res1[9536]);
multi_7x28 multi_7x28_mod_9537(clk,rst,matrix_A[9537],matrix_B[137],mul_res1[9537]);
multi_7x28 multi_7x28_mod_9538(clk,rst,matrix_A[9538],matrix_B[138],mul_res1[9538]);
multi_7x28 multi_7x28_mod_9539(clk,rst,matrix_A[9539],matrix_B[139],mul_res1[9539]);
multi_7x28 multi_7x28_mod_9540(clk,rst,matrix_A[9540],matrix_B[140],mul_res1[9540]);
multi_7x28 multi_7x28_mod_9541(clk,rst,matrix_A[9541],matrix_B[141],mul_res1[9541]);
multi_7x28 multi_7x28_mod_9542(clk,rst,matrix_A[9542],matrix_B[142],mul_res1[9542]);
multi_7x28 multi_7x28_mod_9543(clk,rst,matrix_A[9543],matrix_B[143],mul_res1[9543]);
multi_7x28 multi_7x28_mod_9544(clk,rst,matrix_A[9544],matrix_B[144],mul_res1[9544]);
multi_7x28 multi_7x28_mod_9545(clk,rst,matrix_A[9545],matrix_B[145],mul_res1[9545]);
multi_7x28 multi_7x28_mod_9546(clk,rst,matrix_A[9546],matrix_B[146],mul_res1[9546]);
multi_7x28 multi_7x28_mod_9547(clk,rst,matrix_A[9547],matrix_B[147],mul_res1[9547]);
multi_7x28 multi_7x28_mod_9548(clk,rst,matrix_A[9548],matrix_B[148],mul_res1[9548]);
multi_7x28 multi_7x28_mod_9549(clk,rst,matrix_A[9549],matrix_B[149],mul_res1[9549]);
multi_7x28 multi_7x28_mod_9550(clk,rst,matrix_A[9550],matrix_B[150],mul_res1[9550]);
multi_7x28 multi_7x28_mod_9551(clk,rst,matrix_A[9551],matrix_B[151],mul_res1[9551]);
multi_7x28 multi_7x28_mod_9552(clk,rst,matrix_A[9552],matrix_B[152],mul_res1[9552]);
multi_7x28 multi_7x28_mod_9553(clk,rst,matrix_A[9553],matrix_B[153],mul_res1[9553]);
multi_7x28 multi_7x28_mod_9554(clk,rst,matrix_A[9554],matrix_B[154],mul_res1[9554]);
multi_7x28 multi_7x28_mod_9555(clk,rst,matrix_A[9555],matrix_B[155],mul_res1[9555]);
multi_7x28 multi_7x28_mod_9556(clk,rst,matrix_A[9556],matrix_B[156],mul_res1[9556]);
multi_7x28 multi_7x28_mod_9557(clk,rst,matrix_A[9557],matrix_B[157],mul_res1[9557]);
multi_7x28 multi_7x28_mod_9558(clk,rst,matrix_A[9558],matrix_B[158],mul_res1[9558]);
multi_7x28 multi_7x28_mod_9559(clk,rst,matrix_A[9559],matrix_B[159],mul_res1[9559]);
multi_7x28 multi_7x28_mod_9560(clk,rst,matrix_A[9560],matrix_B[160],mul_res1[9560]);
multi_7x28 multi_7x28_mod_9561(clk,rst,matrix_A[9561],matrix_B[161],mul_res1[9561]);
multi_7x28 multi_7x28_mod_9562(clk,rst,matrix_A[9562],matrix_B[162],mul_res1[9562]);
multi_7x28 multi_7x28_mod_9563(clk,rst,matrix_A[9563],matrix_B[163],mul_res1[9563]);
multi_7x28 multi_7x28_mod_9564(clk,rst,matrix_A[9564],matrix_B[164],mul_res1[9564]);
multi_7x28 multi_7x28_mod_9565(clk,rst,matrix_A[9565],matrix_B[165],mul_res1[9565]);
multi_7x28 multi_7x28_mod_9566(clk,rst,matrix_A[9566],matrix_B[166],mul_res1[9566]);
multi_7x28 multi_7x28_mod_9567(clk,rst,matrix_A[9567],matrix_B[167],mul_res1[9567]);
multi_7x28 multi_7x28_mod_9568(clk,rst,matrix_A[9568],matrix_B[168],mul_res1[9568]);
multi_7x28 multi_7x28_mod_9569(clk,rst,matrix_A[9569],matrix_B[169],mul_res1[9569]);
multi_7x28 multi_7x28_mod_9570(clk,rst,matrix_A[9570],matrix_B[170],mul_res1[9570]);
multi_7x28 multi_7x28_mod_9571(clk,rst,matrix_A[9571],matrix_B[171],mul_res1[9571]);
multi_7x28 multi_7x28_mod_9572(clk,rst,matrix_A[9572],matrix_B[172],mul_res1[9572]);
multi_7x28 multi_7x28_mod_9573(clk,rst,matrix_A[9573],matrix_B[173],mul_res1[9573]);
multi_7x28 multi_7x28_mod_9574(clk,rst,matrix_A[9574],matrix_B[174],mul_res1[9574]);
multi_7x28 multi_7x28_mod_9575(clk,rst,matrix_A[9575],matrix_B[175],mul_res1[9575]);
multi_7x28 multi_7x28_mod_9576(clk,rst,matrix_A[9576],matrix_B[176],mul_res1[9576]);
multi_7x28 multi_7x28_mod_9577(clk,rst,matrix_A[9577],matrix_B[177],mul_res1[9577]);
multi_7x28 multi_7x28_mod_9578(clk,rst,matrix_A[9578],matrix_B[178],mul_res1[9578]);
multi_7x28 multi_7x28_mod_9579(clk,rst,matrix_A[9579],matrix_B[179],mul_res1[9579]);
multi_7x28 multi_7x28_mod_9580(clk,rst,matrix_A[9580],matrix_B[180],mul_res1[9580]);
multi_7x28 multi_7x28_mod_9581(clk,rst,matrix_A[9581],matrix_B[181],mul_res1[9581]);
multi_7x28 multi_7x28_mod_9582(clk,rst,matrix_A[9582],matrix_B[182],mul_res1[9582]);
multi_7x28 multi_7x28_mod_9583(clk,rst,matrix_A[9583],matrix_B[183],mul_res1[9583]);
multi_7x28 multi_7x28_mod_9584(clk,rst,matrix_A[9584],matrix_B[184],mul_res1[9584]);
multi_7x28 multi_7x28_mod_9585(clk,rst,matrix_A[9585],matrix_B[185],mul_res1[9585]);
multi_7x28 multi_7x28_mod_9586(clk,rst,matrix_A[9586],matrix_B[186],mul_res1[9586]);
multi_7x28 multi_7x28_mod_9587(clk,rst,matrix_A[9587],matrix_B[187],mul_res1[9587]);
multi_7x28 multi_7x28_mod_9588(clk,rst,matrix_A[9588],matrix_B[188],mul_res1[9588]);
multi_7x28 multi_7x28_mod_9589(clk,rst,matrix_A[9589],matrix_B[189],mul_res1[9589]);
multi_7x28 multi_7x28_mod_9590(clk,rst,matrix_A[9590],matrix_B[190],mul_res1[9590]);
multi_7x28 multi_7x28_mod_9591(clk,rst,matrix_A[9591],matrix_B[191],mul_res1[9591]);
multi_7x28 multi_7x28_mod_9592(clk,rst,matrix_A[9592],matrix_B[192],mul_res1[9592]);
multi_7x28 multi_7x28_mod_9593(clk,rst,matrix_A[9593],matrix_B[193],mul_res1[9593]);
multi_7x28 multi_7x28_mod_9594(clk,rst,matrix_A[9594],matrix_B[194],mul_res1[9594]);
multi_7x28 multi_7x28_mod_9595(clk,rst,matrix_A[9595],matrix_B[195],mul_res1[9595]);
multi_7x28 multi_7x28_mod_9596(clk,rst,matrix_A[9596],matrix_B[196],mul_res1[9596]);
multi_7x28 multi_7x28_mod_9597(clk,rst,matrix_A[9597],matrix_B[197],mul_res1[9597]);
multi_7x28 multi_7x28_mod_9598(clk,rst,matrix_A[9598],matrix_B[198],mul_res1[9598]);
multi_7x28 multi_7x28_mod_9599(clk,rst,matrix_A[9599],matrix_B[199],mul_res1[9599]);
multi_7x28 multi_7x28_mod_9600(clk,rst,matrix_A[9600],matrix_B[0],mul_res1[9600]);
multi_7x28 multi_7x28_mod_9601(clk,rst,matrix_A[9601],matrix_B[1],mul_res1[9601]);
multi_7x28 multi_7x28_mod_9602(clk,rst,matrix_A[9602],matrix_B[2],mul_res1[9602]);
multi_7x28 multi_7x28_mod_9603(clk,rst,matrix_A[9603],matrix_B[3],mul_res1[9603]);
multi_7x28 multi_7x28_mod_9604(clk,rst,matrix_A[9604],matrix_B[4],mul_res1[9604]);
multi_7x28 multi_7x28_mod_9605(clk,rst,matrix_A[9605],matrix_B[5],mul_res1[9605]);
multi_7x28 multi_7x28_mod_9606(clk,rst,matrix_A[9606],matrix_B[6],mul_res1[9606]);
multi_7x28 multi_7x28_mod_9607(clk,rst,matrix_A[9607],matrix_B[7],mul_res1[9607]);
multi_7x28 multi_7x28_mod_9608(clk,rst,matrix_A[9608],matrix_B[8],mul_res1[9608]);
multi_7x28 multi_7x28_mod_9609(clk,rst,matrix_A[9609],matrix_B[9],mul_res1[9609]);
multi_7x28 multi_7x28_mod_9610(clk,rst,matrix_A[9610],matrix_B[10],mul_res1[9610]);
multi_7x28 multi_7x28_mod_9611(clk,rst,matrix_A[9611],matrix_B[11],mul_res1[9611]);
multi_7x28 multi_7x28_mod_9612(clk,rst,matrix_A[9612],matrix_B[12],mul_res1[9612]);
multi_7x28 multi_7x28_mod_9613(clk,rst,matrix_A[9613],matrix_B[13],mul_res1[9613]);
multi_7x28 multi_7x28_mod_9614(clk,rst,matrix_A[9614],matrix_B[14],mul_res1[9614]);
multi_7x28 multi_7x28_mod_9615(clk,rst,matrix_A[9615],matrix_B[15],mul_res1[9615]);
multi_7x28 multi_7x28_mod_9616(clk,rst,matrix_A[9616],matrix_B[16],mul_res1[9616]);
multi_7x28 multi_7x28_mod_9617(clk,rst,matrix_A[9617],matrix_B[17],mul_res1[9617]);
multi_7x28 multi_7x28_mod_9618(clk,rst,matrix_A[9618],matrix_B[18],mul_res1[9618]);
multi_7x28 multi_7x28_mod_9619(clk,rst,matrix_A[9619],matrix_B[19],mul_res1[9619]);
multi_7x28 multi_7x28_mod_9620(clk,rst,matrix_A[9620],matrix_B[20],mul_res1[9620]);
multi_7x28 multi_7x28_mod_9621(clk,rst,matrix_A[9621],matrix_B[21],mul_res1[9621]);
multi_7x28 multi_7x28_mod_9622(clk,rst,matrix_A[9622],matrix_B[22],mul_res1[9622]);
multi_7x28 multi_7x28_mod_9623(clk,rst,matrix_A[9623],matrix_B[23],mul_res1[9623]);
multi_7x28 multi_7x28_mod_9624(clk,rst,matrix_A[9624],matrix_B[24],mul_res1[9624]);
multi_7x28 multi_7x28_mod_9625(clk,rst,matrix_A[9625],matrix_B[25],mul_res1[9625]);
multi_7x28 multi_7x28_mod_9626(clk,rst,matrix_A[9626],matrix_B[26],mul_res1[9626]);
multi_7x28 multi_7x28_mod_9627(clk,rst,matrix_A[9627],matrix_B[27],mul_res1[9627]);
multi_7x28 multi_7x28_mod_9628(clk,rst,matrix_A[9628],matrix_B[28],mul_res1[9628]);
multi_7x28 multi_7x28_mod_9629(clk,rst,matrix_A[9629],matrix_B[29],mul_res1[9629]);
multi_7x28 multi_7x28_mod_9630(clk,rst,matrix_A[9630],matrix_B[30],mul_res1[9630]);
multi_7x28 multi_7x28_mod_9631(clk,rst,matrix_A[9631],matrix_B[31],mul_res1[9631]);
multi_7x28 multi_7x28_mod_9632(clk,rst,matrix_A[9632],matrix_B[32],mul_res1[9632]);
multi_7x28 multi_7x28_mod_9633(clk,rst,matrix_A[9633],matrix_B[33],mul_res1[9633]);
multi_7x28 multi_7x28_mod_9634(clk,rst,matrix_A[9634],matrix_B[34],mul_res1[9634]);
multi_7x28 multi_7x28_mod_9635(clk,rst,matrix_A[9635],matrix_B[35],mul_res1[9635]);
multi_7x28 multi_7x28_mod_9636(clk,rst,matrix_A[9636],matrix_B[36],mul_res1[9636]);
multi_7x28 multi_7x28_mod_9637(clk,rst,matrix_A[9637],matrix_B[37],mul_res1[9637]);
multi_7x28 multi_7x28_mod_9638(clk,rst,matrix_A[9638],matrix_B[38],mul_res1[9638]);
multi_7x28 multi_7x28_mod_9639(clk,rst,matrix_A[9639],matrix_B[39],mul_res1[9639]);
multi_7x28 multi_7x28_mod_9640(clk,rst,matrix_A[9640],matrix_B[40],mul_res1[9640]);
multi_7x28 multi_7x28_mod_9641(clk,rst,matrix_A[9641],matrix_B[41],mul_res1[9641]);
multi_7x28 multi_7x28_mod_9642(clk,rst,matrix_A[9642],matrix_B[42],mul_res1[9642]);
multi_7x28 multi_7x28_mod_9643(clk,rst,matrix_A[9643],matrix_B[43],mul_res1[9643]);
multi_7x28 multi_7x28_mod_9644(clk,rst,matrix_A[9644],matrix_B[44],mul_res1[9644]);
multi_7x28 multi_7x28_mod_9645(clk,rst,matrix_A[9645],matrix_B[45],mul_res1[9645]);
multi_7x28 multi_7x28_mod_9646(clk,rst,matrix_A[9646],matrix_B[46],mul_res1[9646]);
multi_7x28 multi_7x28_mod_9647(clk,rst,matrix_A[9647],matrix_B[47],mul_res1[9647]);
multi_7x28 multi_7x28_mod_9648(clk,rst,matrix_A[9648],matrix_B[48],mul_res1[9648]);
multi_7x28 multi_7x28_mod_9649(clk,rst,matrix_A[9649],matrix_B[49],mul_res1[9649]);
multi_7x28 multi_7x28_mod_9650(clk,rst,matrix_A[9650],matrix_B[50],mul_res1[9650]);
multi_7x28 multi_7x28_mod_9651(clk,rst,matrix_A[9651],matrix_B[51],mul_res1[9651]);
multi_7x28 multi_7x28_mod_9652(clk,rst,matrix_A[9652],matrix_B[52],mul_res1[9652]);
multi_7x28 multi_7x28_mod_9653(clk,rst,matrix_A[9653],matrix_B[53],mul_res1[9653]);
multi_7x28 multi_7x28_mod_9654(clk,rst,matrix_A[9654],matrix_B[54],mul_res1[9654]);
multi_7x28 multi_7x28_mod_9655(clk,rst,matrix_A[9655],matrix_B[55],mul_res1[9655]);
multi_7x28 multi_7x28_mod_9656(clk,rst,matrix_A[9656],matrix_B[56],mul_res1[9656]);
multi_7x28 multi_7x28_mod_9657(clk,rst,matrix_A[9657],matrix_B[57],mul_res1[9657]);
multi_7x28 multi_7x28_mod_9658(clk,rst,matrix_A[9658],matrix_B[58],mul_res1[9658]);
multi_7x28 multi_7x28_mod_9659(clk,rst,matrix_A[9659],matrix_B[59],mul_res1[9659]);
multi_7x28 multi_7x28_mod_9660(clk,rst,matrix_A[9660],matrix_B[60],mul_res1[9660]);
multi_7x28 multi_7x28_mod_9661(clk,rst,matrix_A[9661],matrix_B[61],mul_res1[9661]);
multi_7x28 multi_7x28_mod_9662(clk,rst,matrix_A[9662],matrix_B[62],mul_res1[9662]);
multi_7x28 multi_7x28_mod_9663(clk,rst,matrix_A[9663],matrix_B[63],mul_res1[9663]);
multi_7x28 multi_7x28_mod_9664(clk,rst,matrix_A[9664],matrix_B[64],mul_res1[9664]);
multi_7x28 multi_7x28_mod_9665(clk,rst,matrix_A[9665],matrix_B[65],mul_res1[9665]);
multi_7x28 multi_7x28_mod_9666(clk,rst,matrix_A[9666],matrix_B[66],mul_res1[9666]);
multi_7x28 multi_7x28_mod_9667(clk,rst,matrix_A[9667],matrix_B[67],mul_res1[9667]);
multi_7x28 multi_7x28_mod_9668(clk,rst,matrix_A[9668],matrix_B[68],mul_res1[9668]);
multi_7x28 multi_7x28_mod_9669(clk,rst,matrix_A[9669],matrix_B[69],mul_res1[9669]);
multi_7x28 multi_7x28_mod_9670(clk,rst,matrix_A[9670],matrix_B[70],mul_res1[9670]);
multi_7x28 multi_7x28_mod_9671(clk,rst,matrix_A[9671],matrix_B[71],mul_res1[9671]);
multi_7x28 multi_7x28_mod_9672(clk,rst,matrix_A[9672],matrix_B[72],mul_res1[9672]);
multi_7x28 multi_7x28_mod_9673(clk,rst,matrix_A[9673],matrix_B[73],mul_res1[9673]);
multi_7x28 multi_7x28_mod_9674(clk,rst,matrix_A[9674],matrix_B[74],mul_res1[9674]);
multi_7x28 multi_7x28_mod_9675(clk,rst,matrix_A[9675],matrix_B[75],mul_res1[9675]);
multi_7x28 multi_7x28_mod_9676(clk,rst,matrix_A[9676],matrix_B[76],mul_res1[9676]);
multi_7x28 multi_7x28_mod_9677(clk,rst,matrix_A[9677],matrix_B[77],mul_res1[9677]);
multi_7x28 multi_7x28_mod_9678(clk,rst,matrix_A[9678],matrix_B[78],mul_res1[9678]);
multi_7x28 multi_7x28_mod_9679(clk,rst,matrix_A[9679],matrix_B[79],mul_res1[9679]);
multi_7x28 multi_7x28_mod_9680(clk,rst,matrix_A[9680],matrix_B[80],mul_res1[9680]);
multi_7x28 multi_7x28_mod_9681(clk,rst,matrix_A[9681],matrix_B[81],mul_res1[9681]);
multi_7x28 multi_7x28_mod_9682(clk,rst,matrix_A[9682],matrix_B[82],mul_res1[9682]);
multi_7x28 multi_7x28_mod_9683(clk,rst,matrix_A[9683],matrix_B[83],mul_res1[9683]);
multi_7x28 multi_7x28_mod_9684(clk,rst,matrix_A[9684],matrix_B[84],mul_res1[9684]);
multi_7x28 multi_7x28_mod_9685(clk,rst,matrix_A[9685],matrix_B[85],mul_res1[9685]);
multi_7x28 multi_7x28_mod_9686(clk,rst,matrix_A[9686],matrix_B[86],mul_res1[9686]);
multi_7x28 multi_7x28_mod_9687(clk,rst,matrix_A[9687],matrix_B[87],mul_res1[9687]);
multi_7x28 multi_7x28_mod_9688(clk,rst,matrix_A[9688],matrix_B[88],mul_res1[9688]);
multi_7x28 multi_7x28_mod_9689(clk,rst,matrix_A[9689],matrix_B[89],mul_res1[9689]);
multi_7x28 multi_7x28_mod_9690(clk,rst,matrix_A[9690],matrix_B[90],mul_res1[9690]);
multi_7x28 multi_7x28_mod_9691(clk,rst,matrix_A[9691],matrix_B[91],mul_res1[9691]);
multi_7x28 multi_7x28_mod_9692(clk,rst,matrix_A[9692],matrix_B[92],mul_res1[9692]);
multi_7x28 multi_7x28_mod_9693(clk,rst,matrix_A[9693],matrix_B[93],mul_res1[9693]);
multi_7x28 multi_7x28_mod_9694(clk,rst,matrix_A[9694],matrix_B[94],mul_res1[9694]);
multi_7x28 multi_7x28_mod_9695(clk,rst,matrix_A[9695],matrix_B[95],mul_res1[9695]);
multi_7x28 multi_7x28_mod_9696(clk,rst,matrix_A[9696],matrix_B[96],mul_res1[9696]);
multi_7x28 multi_7x28_mod_9697(clk,rst,matrix_A[9697],matrix_B[97],mul_res1[9697]);
multi_7x28 multi_7x28_mod_9698(clk,rst,matrix_A[9698],matrix_B[98],mul_res1[9698]);
multi_7x28 multi_7x28_mod_9699(clk,rst,matrix_A[9699],matrix_B[99],mul_res1[9699]);
multi_7x28 multi_7x28_mod_9700(clk,rst,matrix_A[9700],matrix_B[100],mul_res1[9700]);
multi_7x28 multi_7x28_mod_9701(clk,rst,matrix_A[9701],matrix_B[101],mul_res1[9701]);
multi_7x28 multi_7x28_mod_9702(clk,rst,matrix_A[9702],matrix_B[102],mul_res1[9702]);
multi_7x28 multi_7x28_mod_9703(clk,rst,matrix_A[9703],matrix_B[103],mul_res1[9703]);
multi_7x28 multi_7x28_mod_9704(clk,rst,matrix_A[9704],matrix_B[104],mul_res1[9704]);
multi_7x28 multi_7x28_mod_9705(clk,rst,matrix_A[9705],matrix_B[105],mul_res1[9705]);
multi_7x28 multi_7x28_mod_9706(clk,rst,matrix_A[9706],matrix_B[106],mul_res1[9706]);
multi_7x28 multi_7x28_mod_9707(clk,rst,matrix_A[9707],matrix_B[107],mul_res1[9707]);
multi_7x28 multi_7x28_mod_9708(clk,rst,matrix_A[9708],matrix_B[108],mul_res1[9708]);
multi_7x28 multi_7x28_mod_9709(clk,rst,matrix_A[9709],matrix_B[109],mul_res1[9709]);
multi_7x28 multi_7x28_mod_9710(clk,rst,matrix_A[9710],matrix_B[110],mul_res1[9710]);
multi_7x28 multi_7x28_mod_9711(clk,rst,matrix_A[9711],matrix_B[111],mul_res1[9711]);
multi_7x28 multi_7x28_mod_9712(clk,rst,matrix_A[9712],matrix_B[112],mul_res1[9712]);
multi_7x28 multi_7x28_mod_9713(clk,rst,matrix_A[9713],matrix_B[113],mul_res1[9713]);
multi_7x28 multi_7x28_mod_9714(clk,rst,matrix_A[9714],matrix_B[114],mul_res1[9714]);
multi_7x28 multi_7x28_mod_9715(clk,rst,matrix_A[9715],matrix_B[115],mul_res1[9715]);
multi_7x28 multi_7x28_mod_9716(clk,rst,matrix_A[9716],matrix_B[116],mul_res1[9716]);
multi_7x28 multi_7x28_mod_9717(clk,rst,matrix_A[9717],matrix_B[117],mul_res1[9717]);
multi_7x28 multi_7x28_mod_9718(clk,rst,matrix_A[9718],matrix_B[118],mul_res1[9718]);
multi_7x28 multi_7x28_mod_9719(clk,rst,matrix_A[9719],matrix_B[119],mul_res1[9719]);
multi_7x28 multi_7x28_mod_9720(clk,rst,matrix_A[9720],matrix_B[120],mul_res1[9720]);
multi_7x28 multi_7x28_mod_9721(clk,rst,matrix_A[9721],matrix_B[121],mul_res1[9721]);
multi_7x28 multi_7x28_mod_9722(clk,rst,matrix_A[9722],matrix_B[122],mul_res1[9722]);
multi_7x28 multi_7x28_mod_9723(clk,rst,matrix_A[9723],matrix_B[123],mul_res1[9723]);
multi_7x28 multi_7x28_mod_9724(clk,rst,matrix_A[9724],matrix_B[124],mul_res1[9724]);
multi_7x28 multi_7x28_mod_9725(clk,rst,matrix_A[9725],matrix_B[125],mul_res1[9725]);
multi_7x28 multi_7x28_mod_9726(clk,rst,matrix_A[9726],matrix_B[126],mul_res1[9726]);
multi_7x28 multi_7x28_mod_9727(clk,rst,matrix_A[9727],matrix_B[127],mul_res1[9727]);
multi_7x28 multi_7x28_mod_9728(clk,rst,matrix_A[9728],matrix_B[128],mul_res1[9728]);
multi_7x28 multi_7x28_mod_9729(clk,rst,matrix_A[9729],matrix_B[129],mul_res1[9729]);
multi_7x28 multi_7x28_mod_9730(clk,rst,matrix_A[9730],matrix_B[130],mul_res1[9730]);
multi_7x28 multi_7x28_mod_9731(clk,rst,matrix_A[9731],matrix_B[131],mul_res1[9731]);
multi_7x28 multi_7x28_mod_9732(clk,rst,matrix_A[9732],matrix_B[132],mul_res1[9732]);
multi_7x28 multi_7x28_mod_9733(clk,rst,matrix_A[9733],matrix_B[133],mul_res1[9733]);
multi_7x28 multi_7x28_mod_9734(clk,rst,matrix_A[9734],matrix_B[134],mul_res1[9734]);
multi_7x28 multi_7x28_mod_9735(clk,rst,matrix_A[9735],matrix_B[135],mul_res1[9735]);
multi_7x28 multi_7x28_mod_9736(clk,rst,matrix_A[9736],matrix_B[136],mul_res1[9736]);
multi_7x28 multi_7x28_mod_9737(clk,rst,matrix_A[9737],matrix_B[137],mul_res1[9737]);
multi_7x28 multi_7x28_mod_9738(clk,rst,matrix_A[9738],matrix_B[138],mul_res1[9738]);
multi_7x28 multi_7x28_mod_9739(clk,rst,matrix_A[9739],matrix_B[139],mul_res1[9739]);
multi_7x28 multi_7x28_mod_9740(clk,rst,matrix_A[9740],matrix_B[140],mul_res1[9740]);
multi_7x28 multi_7x28_mod_9741(clk,rst,matrix_A[9741],matrix_B[141],mul_res1[9741]);
multi_7x28 multi_7x28_mod_9742(clk,rst,matrix_A[9742],matrix_B[142],mul_res1[9742]);
multi_7x28 multi_7x28_mod_9743(clk,rst,matrix_A[9743],matrix_B[143],mul_res1[9743]);
multi_7x28 multi_7x28_mod_9744(clk,rst,matrix_A[9744],matrix_B[144],mul_res1[9744]);
multi_7x28 multi_7x28_mod_9745(clk,rst,matrix_A[9745],matrix_B[145],mul_res1[9745]);
multi_7x28 multi_7x28_mod_9746(clk,rst,matrix_A[9746],matrix_B[146],mul_res1[9746]);
multi_7x28 multi_7x28_mod_9747(clk,rst,matrix_A[9747],matrix_B[147],mul_res1[9747]);
multi_7x28 multi_7x28_mod_9748(clk,rst,matrix_A[9748],matrix_B[148],mul_res1[9748]);
multi_7x28 multi_7x28_mod_9749(clk,rst,matrix_A[9749],matrix_B[149],mul_res1[9749]);
multi_7x28 multi_7x28_mod_9750(clk,rst,matrix_A[9750],matrix_B[150],mul_res1[9750]);
multi_7x28 multi_7x28_mod_9751(clk,rst,matrix_A[9751],matrix_B[151],mul_res1[9751]);
multi_7x28 multi_7x28_mod_9752(clk,rst,matrix_A[9752],matrix_B[152],mul_res1[9752]);
multi_7x28 multi_7x28_mod_9753(clk,rst,matrix_A[9753],matrix_B[153],mul_res1[9753]);
multi_7x28 multi_7x28_mod_9754(clk,rst,matrix_A[9754],matrix_B[154],mul_res1[9754]);
multi_7x28 multi_7x28_mod_9755(clk,rst,matrix_A[9755],matrix_B[155],mul_res1[9755]);
multi_7x28 multi_7x28_mod_9756(clk,rst,matrix_A[9756],matrix_B[156],mul_res1[9756]);
multi_7x28 multi_7x28_mod_9757(clk,rst,matrix_A[9757],matrix_B[157],mul_res1[9757]);
multi_7x28 multi_7x28_mod_9758(clk,rst,matrix_A[9758],matrix_B[158],mul_res1[9758]);
multi_7x28 multi_7x28_mod_9759(clk,rst,matrix_A[9759],matrix_B[159],mul_res1[9759]);
multi_7x28 multi_7x28_mod_9760(clk,rst,matrix_A[9760],matrix_B[160],mul_res1[9760]);
multi_7x28 multi_7x28_mod_9761(clk,rst,matrix_A[9761],matrix_B[161],mul_res1[9761]);
multi_7x28 multi_7x28_mod_9762(clk,rst,matrix_A[9762],matrix_B[162],mul_res1[9762]);
multi_7x28 multi_7x28_mod_9763(clk,rst,matrix_A[9763],matrix_B[163],mul_res1[9763]);
multi_7x28 multi_7x28_mod_9764(clk,rst,matrix_A[9764],matrix_B[164],mul_res1[9764]);
multi_7x28 multi_7x28_mod_9765(clk,rst,matrix_A[9765],matrix_B[165],mul_res1[9765]);
multi_7x28 multi_7x28_mod_9766(clk,rst,matrix_A[9766],matrix_B[166],mul_res1[9766]);
multi_7x28 multi_7x28_mod_9767(clk,rst,matrix_A[9767],matrix_B[167],mul_res1[9767]);
multi_7x28 multi_7x28_mod_9768(clk,rst,matrix_A[9768],matrix_B[168],mul_res1[9768]);
multi_7x28 multi_7x28_mod_9769(clk,rst,matrix_A[9769],matrix_B[169],mul_res1[9769]);
multi_7x28 multi_7x28_mod_9770(clk,rst,matrix_A[9770],matrix_B[170],mul_res1[9770]);
multi_7x28 multi_7x28_mod_9771(clk,rst,matrix_A[9771],matrix_B[171],mul_res1[9771]);
multi_7x28 multi_7x28_mod_9772(clk,rst,matrix_A[9772],matrix_B[172],mul_res1[9772]);
multi_7x28 multi_7x28_mod_9773(clk,rst,matrix_A[9773],matrix_B[173],mul_res1[9773]);
multi_7x28 multi_7x28_mod_9774(clk,rst,matrix_A[9774],matrix_B[174],mul_res1[9774]);
multi_7x28 multi_7x28_mod_9775(clk,rst,matrix_A[9775],matrix_B[175],mul_res1[9775]);
multi_7x28 multi_7x28_mod_9776(clk,rst,matrix_A[9776],matrix_B[176],mul_res1[9776]);
multi_7x28 multi_7x28_mod_9777(clk,rst,matrix_A[9777],matrix_B[177],mul_res1[9777]);
multi_7x28 multi_7x28_mod_9778(clk,rst,matrix_A[9778],matrix_B[178],mul_res1[9778]);
multi_7x28 multi_7x28_mod_9779(clk,rst,matrix_A[9779],matrix_B[179],mul_res1[9779]);
multi_7x28 multi_7x28_mod_9780(clk,rst,matrix_A[9780],matrix_B[180],mul_res1[9780]);
multi_7x28 multi_7x28_mod_9781(clk,rst,matrix_A[9781],matrix_B[181],mul_res1[9781]);
multi_7x28 multi_7x28_mod_9782(clk,rst,matrix_A[9782],matrix_B[182],mul_res1[9782]);
multi_7x28 multi_7x28_mod_9783(clk,rst,matrix_A[9783],matrix_B[183],mul_res1[9783]);
multi_7x28 multi_7x28_mod_9784(clk,rst,matrix_A[9784],matrix_B[184],mul_res1[9784]);
multi_7x28 multi_7x28_mod_9785(clk,rst,matrix_A[9785],matrix_B[185],mul_res1[9785]);
multi_7x28 multi_7x28_mod_9786(clk,rst,matrix_A[9786],matrix_B[186],mul_res1[9786]);
multi_7x28 multi_7x28_mod_9787(clk,rst,matrix_A[9787],matrix_B[187],mul_res1[9787]);
multi_7x28 multi_7x28_mod_9788(clk,rst,matrix_A[9788],matrix_B[188],mul_res1[9788]);
multi_7x28 multi_7x28_mod_9789(clk,rst,matrix_A[9789],matrix_B[189],mul_res1[9789]);
multi_7x28 multi_7x28_mod_9790(clk,rst,matrix_A[9790],matrix_B[190],mul_res1[9790]);
multi_7x28 multi_7x28_mod_9791(clk,rst,matrix_A[9791],matrix_B[191],mul_res1[9791]);
multi_7x28 multi_7x28_mod_9792(clk,rst,matrix_A[9792],matrix_B[192],mul_res1[9792]);
multi_7x28 multi_7x28_mod_9793(clk,rst,matrix_A[9793],matrix_B[193],mul_res1[9793]);
multi_7x28 multi_7x28_mod_9794(clk,rst,matrix_A[9794],matrix_B[194],mul_res1[9794]);
multi_7x28 multi_7x28_mod_9795(clk,rst,matrix_A[9795],matrix_B[195],mul_res1[9795]);
multi_7x28 multi_7x28_mod_9796(clk,rst,matrix_A[9796],matrix_B[196],mul_res1[9796]);
multi_7x28 multi_7x28_mod_9797(clk,rst,matrix_A[9797],matrix_B[197],mul_res1[9797]);
multi_7x28 multi_7x28_mod_9798(clk,rst,matrix_A[9798],matrix_B[198],mul_res1[9798]);
multi_7x28 multi_7x28_mod_9799(clk,rst,matrix_A[9799],matrix_B[199],mul_res1[9799]);
multi_7x28 multi_7x28_mod_9800(clk,rst,matrix_A[9800],matrix_B[0],mul_res1[9800]);
multi_7x28 multi_7x28_mod_9801(clk,rst,matrix_A[9801],matrix_B[1],mul_res1[9801]);
multi_7x28 multi_7x28_mod_9802(clk,rst,matrix_A[9802],matrix_B[2],mul_res1[9802]);
multi_7x28 multi_7x28_mod_9803(clk,rst,matrix_A[9803],matrix_B[3],mul_res1[9803]);
multi_7x28 multi_7x28_mod_9804(clk,rst,matrix_A[9804],matrix_B[4],mul_res1[9804]);
multi_7x28 multi_7x28_mod_9805(clk,rst,matrix_A[9805],matrix_B[5],mul_res1[9805]);
multi_7x28 multi_7x28_mod_9806(clk,rst,matrix_A[9806],matrix_B[6],mul_res1[9806]);
multi_7x28 multi_7x28_mod_9807(clk,rst,matrix_A[9807],matrix_B[7],mul_res1[9807]);
multi_7x28 multi_7x28_mod_9808(clk,rst,matrix_A[9808],matrix_B[8],mul_res1[9808]);
multi_7x28 multi_7x28_mod_9809(clk,rst,matrix_A[9809],matrix_B[9],mul_res1[9809]);
multi_7x28 multi_7x28_mod_9810(clk,rst,matrix_A[9810],matrix_B[10],mul_res1[9810]);
multi_7x28 multi_7x28_mod_9811(clk,rst,matrix_A[9811],matrix_B[11],mul_res1[9811]);
multi_7x28 multi_7x28_mod_9812(clk,rst,matrix_A[9812],matrix_B[12],mul_res1[9812]);
multi_7x28 multi_7x28_mod_9813(clk,rst,matrix_A[9813],matrix_B[13],mul_res1[9813]);
multi_7x28 multi_7x28_mod_9814(clk,rst,matrix_A[9814],matrix_B[14],mul_res1[9814]);
multi_7x28 multi_7x28_mod_9815(clk,rst,matrix_A[9815],matrix_B[15],mul_res1[9815]);
multi_7x28 multi_7x28_mod_9816(clk,rst,matrix_A[9816],matrix_B[16],mul_res1[9816]);
multi_7x28 multi_7x28_mod_9817(clk,rst,matrix_A[9817],matrix_B[17],mul_res1[9817]);
multi_7x28 multi_7x28_mod_9818(clk,rst,matrix_A[9818],matrix_B[18],mul_res1[9818]);
multi_7x28 multi_7x28_mod_9819(clk,rst,matrix_A[9819],matrix_B[19],mul_res1[9819]);
multi_7x28 multi_7x28_mod_9820(clk,rst,matrix_A[9820],matrix_B[20],mul_res1[9820]);
multi_7x28 multi_7x28_mod_9821(clk,rst,matrix_A[9821],matrix_B[21],mul_res1[9821]);
multi_7x28 multi_7x28_mod_9822(clk,rst,matrix_A[9822],matrix_B[22],mul_res1[9822]);
multi_7x28 multi_7x28_mod_9823(clk,rst,matrix_A[9823],matrix_B[23],mul_res1[9823]);
multi_7x28 multi_7x28_mod_9824(clk,rst,matrix_A[9824],matrix_B[24],mul_res1[9824]);
multi_7x28 multi_7x28_mod_9825(clk,rst,matrix_A[9825],matrix_B[25],mul_res1[9825]);
multi_7x28 multi_7x28_mod_9826(clk,rst,matrix_A[9826],matrix_B[26],mul_res1[9826]);
multi_7x28 multi_7x28_mod_9827(clk,rst,matrix_A[9827],matrix_B[27],mul_res1[9827]);
multi_7x28 multi_7x28_mod_9828(clk,rst,matrix_A[9828],matrix_B[28],mul_res1[9828]);
multi_7x28 multi_7x28_mod_9829(clk,rst,matrix_A[9829],matrix_B[29],mul_res1[9829]);
multi_7x28 multi_7x28_mod_9830(clk,rst,matrix_A[9830],matrix_B[30],mul_res1[9830]);
multi_7x28 multi_7x28_mod_9831(clk,rst,matrix_A[9831],matrix_B[31],mul_res1[9831]);
multi_7x28 multi_7x28_mod_9832(clk,rst,matrix_A[9832],matrix_B[32],mul_res1[9832]);
multi_7x28 multi_7x28_mod_9833(clk,rst,matrix_A[9833],matrix_B[33],mul_res1[9833]);
multi_7x28 multi_7x28_mod_9834(clk,rst,matrix_A[9834],matrix_B[34],mul_res1[9834]);
multi_7x28 multi_7x28_mod_9835(clk,rst,matrix_A[9835],matrix_B[35],mul_res1[9835]);
multi_7x28 multi_7x28_mod_9836(clk,rst,matrix_A[9836],matrix_B[36],mul_res1[9836]);
multi_7x28 multi_7x28_mod_9837(clk,rst,matrix_A[9837],matrix_B[37],mul_res1[9837]);
multi_7x28 multi_7x28_mod_9838(clk,rst,matrix_A[9838],matrix_B[38],mul_res1[9838]);
multi_7x28 multi_7x28_mod_9839(clk,rst,matrix_A[9839],matrix_B[39],mul_res1[9839]);
multi_7x28 multi_7x28_mod_9840(clk,rst,matrix_A[9840],matrix_B[40],mul_res1[9840]);
multi_7x28 multi_7x28_mod_9841(clk,rst,matrix_A[9841],matrix_B[41],mul_res1[9841]);
multi_7x28 multi_7x28_mod_9842(clk,rst,matrix_A[9842],matrix_B[42],mul_res1[9842]);
multi_7x28 multi_7x28_mod_9843(clk,rst,matrix_A[9843],matrix_B[43],mul_res1[9843]);
multi_7x28 multi_7x28_mod_9844(clk,rst,matrix_A[9844],matrix_B[44],mul_res1[9844]);
multi_7x28 multi_7x28_mod_9845(clk,rst,matrix_A[9845],matrix_B[45],mul_res1[9845]);
multi_7x28 multi_7x28_mod_9846(clk,rst,matrix_A[9846],matrix_B[46],mul_res1[9846]);
multi_7x28 multi_7x28_mod_9847(clk,rst,matrix_A[9847],matrix_B[47],mul_res1[9847]);
multi_7x28 multi_7x28_mod_9848(clk,rst,matrix_A[9848],matrix_B[48],mul_res1[9848]);
multi_7x28 multi_7x28_mod_9849(clk,rst,matrix_A[9849],matrix_B[49],mul_res1[9849]);
multi_7x28 multi_7x28_mod_9850(clk,rst,matrix_A[9850],matrix_B[50],mul_res1[9850]);
multi_7x28 multi_7x28_mod_9851(clk,rst,matrix_A[9851],matrix_B[51],mul_res1[9851]);
multi_7x28 multi_7x28_mod_9852(clk,rst,matrix_A[9852],matrix_B[52],mul_res1[9852]);
multi_7x28 multi_7x28_mod_9853(clk,rst,matrix_A[9853],matrix_B[53],mul_res1[9853]);
multi_7x28 multi_7x28_mod_9854(clk,rst,matrix_A[9854],matrix_B[54],mul_res1[9854]);
multi_7x28 multi_7x28_mod_9855(clk,rst,matrix_A[9855],matrix_B[55],mul_res1[9855]);
multi_7x28 multi_7x28_mod_9856(clk,rst,matrix_A[9856],matrix_B[56],mul_res1[9856]);
multi_7x28 multi_7x28_mod_9857(clk,rst,matrix_A[9857],matrix_B[57],mul_res1[9857]);
multi_7x28 multi_7x28_mod_9858(clk,rst,matrix_A[9858],matrix_B[58],mul_res1[9858]);
multi_7x28 multi_7x28_mod_9859(clk,rst,matrix_A[9859],matrix_B[59],mul_res1[9859]);
multi_7x28 multi_7x28_mod_9860(clk,rst,matrix_A[9860],matrix_B[60],mul_res1[9860]);
multi_7x28 multi_7x28_mod_9861(clk,rst,matrix_A[9861],matrix_B[61],mul_res1[9861]);
multi_7x28 multi_7x28_mod_9862(clk,rst,matrix_A[9862],matrix_B[62],mul_res1[9862]);
multi_7x28 multi_7x28_mod_9863(clk,rst,matrix_A[9863],matrix_B[63],mul_res1[9863]);
multi_7x28 multi_7x28_mod_9864(clk,rst,matrix_A[9864],matrix_B[64],mul_res1[9864]);
multi_7x28 multi_7x28_mod_9865(clk,rst,matrix_A[9865],matrix_B[65],mul_res1[9865]);
multi_7x28 multi_7x28_mod_9866(clk,rst,matrix_A[9866],matrix_B[66],mul_res1[9866]);
multi_7x28 multi_7x28_mod_9867(clk,rst,matrix_A[9867],matrix_B[67],mul_res1[9867]);
multi_7x28 multi_7x28_mod_9868(clk,rst,matrix_A[9868],matrix_B[68],mul_res1[9868]);
multi_7x28 multi_7x28_mod_9869(clk,rst,matrix_A[9869],matrix_B[69],mul_res1[9869]);
multi_7x28 multi_7x28_mod_9870(clk,rst,matrix_A[9870],matrix_B[70],mul_res1[9870]);
multi_7x28 multi_7x28_mod_9871(clk,rst,matrix_A[9871],matrix_B[71],mul_res1[9871]);
multi_7x28 multi_7x28_mod_9872(clk,rst,matrix_A[9872],matrix_B[72],mul_res1[9872]);
multi_7x28 multi_7x28_mod_9873(clk,rst,matrix_A[9873],matrix_B[73],mul_res1[9873]);
multi_7x28 multi_7x28_mod_9874(clk,rst,matrix_A[9874],matrix_B[74],mul_res1[9874]);
multi_7x28 multi_7x28_mod_9875(clk,rst,matrix_A[9875],matrix_B[75],mul_res1[9875]);
multi_7x28 multi_7x28_mod_9876(clk,rst,matrix_A[9876],matrix_B[76],mul_res1[9876]);
multi_7x28 multi_7x28_mod_9877(clk,rst,matrix_A[9877],matrix_B[77],mul_res1[9877]);
multi_7x28 multi_7x28_mod_9878(clk,rst,matrix_A[9878],matrix_B[78],mul_res1[9878]);
multi_7x28 multi_7x28_mod_9879(clk,rst,matrix_A[9879],matrix_B[79],mul_res1[9879]);
multi_7x28 multi_7x28_mod_9880(clk,rst,matrix_A[9880],matrix_B[80],mul_res1[9880]);
multi_7x28 multi_7x28_mod_9881(clk,rst,matrix_A[9881],matrix_B[81],mul_res1[9881]);
multi_7x28 multi_7x28_mod_9882(clk,rst,matrix_A[9882],matrix_B[82],mul_res1[9882]);
multi_7x28 multi_7x28_mod_9883(clk,rst,matrix_A[9883],matrix_B[83],mul_res1[9883]);
multi_7x28 multi_7x28_mod_9884(clk,rst,matrix_A[9884],matrix_B[84],mul_res1[9884]);
multi_7x28 multi_7x28_mod_9885(clk,rst,matrix_A[9885],matrix_B[85],mul_res1[9885]);
multi_7x28 multi_7x28_mod_9886(clk,rst,matrix_A[9886],matrix_B[86],mul_res1[9886]);
multi_7x28 multi_7x28_mod_9887(clk,rst,matrix_A[9887],matrix_B[87],mul_res1[9887]);
multi_7x28 multi_7x28_mod_9888(clk,rst,matrix_A[9888],matrix_B[88],mul_res1[9888]);
multi_7x28 multi_7x28_mod_9889(clk,rst,matrix_A[9889],matrix_B[89],mul_res1[9889]);
multi_7x28 multi_7x28_mod_9890(clk,rst,matrix_A[9890],matrix_B[90],mul_res1[9890]);
multi_7x28 multi_7x28_mod_9891(clk,rst,matrix_A[9891],matrix_B[91],mul_res1[9891]);
multi_7x28 multi_7x28_mod_9892(clk,rst,matrix_A[9892],matrix_B[92],mul_res1[9892]);
multi_7x28 multi_7x28_mod_9893(clk,rst,matrix_A[9893],matrix_B[93],mul_res1[9893]);
multi_7x28 multi_7x28_mod_9894(clk,rst,matrix_A[9894],matrix_B[94],mul_res1[9894]);
multi_7x28 multi_7x28_mod_9895(clk,rst,matrix_A[9895],matrix_B[95],mul_res1[9895]);
multi_7x28 multi_7x28_mod_9896(clk,rst,matrix_A[9896],matrix_B[96],mul_res1[9896]);
multi_7x28 multi_7x28_mod_9897(clk,rst,matrix_A[9897],matrix_B[97],mul_res1[9897]);
multi_7x28 multi_7x28_mod_9898(clk,rst,matrix_A[9898],matrix_B[98],mul_res1[9898]);
multi_7x28 multi_7x28_mod_9899(clk,rst,matrix_A[9899],matrix_B[99],mul_res1[9899]);
multi_7x28 multi_7x28_mod_9900(clk,rst,matrix_A[9900],matrix_B[100],mul_res1[9900]);
multi_7x28 multi_7x28_mod_9901(clk,rst,matrix_A[9901],matrix_B[101],mul_res1[9901]);
multi_7x28 multi_7x28_mod_9902(clk,rst,matrix_A[9902],matrix_B[102],mul_res1[9902]);
multi_7x28 multi_7x28_mod_9903(clk,rst,matrix_A[9903],matrix_B[103],mul_res1[9903]);
multi_7x28 multi_7x28_mod_9904(clk,rst,matrix_A[9904],matrix_B[104],mul_res1[9904]);
multi_7x28 multi_7x28_mod_9905(clk,rst,matrix_A[9905],matrix_B[105],mul_res1[9905]);
multi_7x28 multi_7x28_mod_9906(clk,rst,matrix_A[9906],matrix_B[106],mul_res1[9906]);
multi_7x28 multi_7x28_mod_9907(clk,rst,matrix_A[9907],matrix_B[107],mul_res1[9907]);
multi_7x28 multi_7x28_mod_9908(clk,rst,matrix_A[9908],matrix_B[108],mul_res1[9908]);
multi_7x28 multi_7x28_mod_9909(clk,rst,matrix_A[9909],matrix_B[109],mul_res1[9909]);
multi_7x28 multi_7x28_mod_9910(clk,rst,matrix_A[9910],matrix_B[110],mul_res1[9910]);
multi_7x28 multi_7x28_mod_9911(clk,rst,matrix_A[9911],matrix_B[111],mul_res1[9911]);
multi_7x28 multi_7x28_mod_9912(clk,rst,matrix_A[9912],matrix_B[112],mul_res1[9912]);
multi_7x28 multi_7x28_mod_9913(clk,rst,matrix_A[9913],matrix_B[113],mul_res1[9913]);
multi_7x28 multi_7x28_mod_9914(clk,rst,matrix_A[9914],matrix_B[114],mul_res1[9914]);
multi_7x28 multi_7x28_mod_9915(clk,rst,matrix_A[9915],matrix_B[115],mul_res1[9915]);
multi_7x28 multi_7x28_mod_9916(clk,rst,matrix_A[9916],matrix_B[116],mul_res1[9916]);
multi_7x28 multi_7x28_mod_9917(clk,rst,matrix_A[9917],matrix_B[117],mul_res1[9917]);
multi_7x28 multi_7x28_mod_9918(clk,rst,matrix_A[9918],matrix_B[118],mul_res1[9918]);
multi_7x28 multi_7x28_mod_9919(clk,rst,matrix_A[9919],matrix_B[119],mul_res1[9919]);
multi_7x28 multi_7x28_mod_9920(clk,rst,matrix_A[9920],matrix_B[120],mul_res1[9920]);
multi_7x28 multi_7x28_mod_9921(clk,rst,matrix_A[9921],matrix_B[121],mul_res1[9921]);
multi_7x28 multi_7x28_mod_9922(clk,rst,matrix_A[9922],matrix_B[122],mul_res1[9922]);
multi_7x28 multi_7x28_mod_9923(clk,rst,matrix_A[9923],matrix_B[123],mul_res1[9923]);
multi_7x28 multi_7x28_mod_9924(clk,rst,matrix_A[9924],matrix_B[124],mul_res1[9924]);
multi_7x28 multi_7x28_mod_9925(clk,rst,matrix_A[9925],matrix_B[125],mul_res1[9925]);
multi_7x28 multi_7x28_mod_9926(clk,rst,matrix_A[9926],matrix_B[126],mul_res1[9926]);
multi_7x28 multi_7x28_mod_9927(clk,rst,matrix_A[9927],matrix_B[127],mul_res1[9927]);
multi_7x28 multi_7x28_mod_9928(clk,rst,matrix_A[9928],matrix_B[128],mul_res1[9928]);
multi_7x28 multi_7x28_mod_9929(clk,rst,matrix_A[9929],matrix_B[129],mul_res1[9929]);
multi_7x28 multi_7x28_mod_9930(clk,rst,matrix_A[9930],matrix_B[130],mul_res1[9930]);
multi_7x28 multi_7x28_mod_9931(clk,rst,matrix_A[9931],matrix_B[131],mul_res1[9931]);
multi_7x28 multi_7x28_mod_9932(clk,rst,matrix_A[9932],matrix_B[132],mul_res1[9932]);
multi_7x28 multi_7x28_mod_9933(clk,rst,matrix_A[9933],matrix_B[133],mul_res1[9933]);
multi_7x28 multi_7x28_mod_9934(clk,rst,matrix_A[9934],matrix_B[134],mul_res1[9934]);
multi_7x28 multi_7x28_mod_9935(clk,rst,matrix_A[9935],matrix_B[135],mul_res1[9935]);
multi_7x28 multi_7x28_mod_9936(clk,rst,matrix_A[9936],matrix_B[136],mul_res1[9936]);
multi_7x28 multi_7x28_mod_9937(clk,rst,matrix_A[9937],matrix_B[137],mul_res1[9937]);
multi_7x28 multi_7x28_mod_9938(clk,rst,matrix_A[9938],matrix_B[138],mul_res1[9938]);
multi_7x28 multi_7x28_mod_9939(clk,rst,matrix_A[9939],matrix_B[139],mul_res1[9939]);
multi_7x28 multi_7x28_mod_9940(clk,rst,matrix_A[9940],matrix_B[140],mul_res1[9940]);
multi_7x28 multi_7x28_mod_9941(clk,rst,matrix_A[9941],matrix_B[141],mul_res1[9941]);
multi_7x28 multi_7x28_mod_9942(clk,rst,matrix_A[9942],matrix_B[142],mul_res1[9942]);
multi_7x28 multi_7x28_mod_9943(clk,rst,matrix_A[9943],matrix_B[143],mul_res1[9943]);
multi_7x28 multi_7x28_mod_9944(clk,rst,matrix_A[9944],matrix_B[144],mul_res1[9944]);
multi_7x28 multi_7x28_mod_9945(clk,rst,matrix_A[9945],matrix_B[145],mul_res1[9945]);
multi_7x28 multi_7x28_mod_9946(clk,rst,matrix_A[9946],matrix_B[146],mul_res1[9946]);
multi_7x28 multi_7x28_mod_9947(clk,rst,matrix_A[9947],matrix_B[147],mul_res1[9947]);
multi_7x28 multi_7x28_mod_9948(clk,rst,matrix_A[9948],matrix_B[148],mul_res1[9948]);
multi_7x28 multi_7x28_mod_9949(clk,rst,matrix_A[9949],matrix_B[149],mul_res1[9949]);
multi_7x28 multi_7x28_mod_9950(clk,rst,matrix_A[9950],matrix_B[150],mul_res1[9950]);
multi_7x28 multi_7x28_mod_9951(clk,rst,matrix_A[9951],matrix_B[151],mul_res1[9951]);
multi_7x28 multi_7x28_mod_9952(clk,rst,matrix_A[9952],matrix_B[152],mul_res1[9952]);
multi_7x28 multi_7x28_mod_9953(clk,rst,matrix_A[9953],matrix_B[153],mul_res1[9953]);
multi_7x28 multi_7x28_mod_9954(clk,rst,matrix_A[9954],matrix_B[154],mul_res1[9954]);
multi_7x28 multi_7x28_mod_9955(clk,rst,matrix_A[9955],matrix_B[155],mul_res1[9955]);
multi_7x28 multi_7x28_mod_9956(clk,rst,matrix_A[9956],matrix_B[156],mul_res1[9956]);
multi_7x28 multi_7x28_mod_9957(clk,rst,matrix_A[9957],matrix_B[157],mul_res1[9957]);
multi_7x28 multi_7x28_mod_9958(clk,rst,matrix_A[9958],matrix_B[158],mul_res1[9958]);
multi_7x28 multi_7x28_mod_9959(clk,rst,matrix_A[9959],matrix_B[159],mul_res1[9959]);
multi_7x28 multi_7x28_mod_9960(clk,rst,matrix_A[9960],matrix_B[160],mul_res1[9960]);
multi_7x28 multi_7x28_mod_9961(clk,rst,matrix_A[9961],matrix_B[161],mul_res1[9961]);
multi_7x28 multi_7x28_mod_9962(clk,rst,matrix_A[9962],matrix_B[162],mul_res1[9962]);
multi_7x28 multi_7x28_mod_9963(clk,rst,matrix_A[9963],matrix_B[163],mul_res1[9963]);
multi_7x28 multi_7x28_mod_9964(clk,rst,matrix_A[9964],matrix_B[164],mul_res1[9964]);
multi_7x28 multi_7x28_mod_9965(clk,rst,matrix_A[9965],matrix_B[165],mul_res1[9965]);
multi_7x28 multi_7x28_mod_9966(clk,rst,matrix_A[9966],matrix_B[166],mul_res1[9966]);
multi_7x28 multi_7x28_mod_9967(clk,rst,matrix_A[9967],matrix_B[167],mul_res1[9967]);
multi_7x28 multi_7x28_mod_9968(clk,rst,matrix_A[9968],matrix_B[168],mul_res1[9968]);
multi_7x28 multi_7x28_mod_9969(clk,rst,matrix_A[9969],matrix_B[169],mul_res1[9969]);
multi_7x28 multi_7x28_mod_9970(clk,rst,matrix_A[9970],matrix_B[170],mul_res1[9970]);
multi_7x28 multi_7x28_mod_9971(clk,rst,matrix_A[9971],matrix_B[171],mul_res1[9971]);
multi_7x28 multi_7x28_mod_9972(clk,rst,matrix_A[9972],matrix_B[172],mul_res1[9972]);
multi_7x28 multi_7x28_mod_9973(clk,rst,matrix_A[9973],matrix_B[173],mul_res1[9973]);
multi_7x28 multi_7x28_mod_9974(clk,rst,matrix_A[9974],matrix_B[174],mul_res1[9974]);
multi_7x28 multi_7x28_mod_9975(clk,rst,matrix_A[9975],matrix_B[175],mul_res1[9975]);
multi_7x28 multi_7x28_mod_9976(clk,rst,matrix_A[9976],matrix_B[176],mul_res1[9976]);
multi_7x28 multi_7x28_mod_9977(clk,rst,matrix_A[9977],matrix_B[177],mul_res1[9977]);
multi_7x28 multi_7x28_mod_9978(clk,rst,matrix_A[9978],matrix_B[178],mul_res1[9978]);
multi_7x28 multi_7x28_mod_9979(clk,rst,matrix_A[9979],matrix_B[179],mul_res1[9979]);
multi_7x28 multi_7x28_mod_9980(clk,rst,matrix_A[9980],matrix_B[180],mul_res1[9980]);
multi_7x28 multi_7x28_mod_9981(clk,rst,matrix_A[9981],matrix_B[181],mul_res1[9981]);
multi_7x28 multi_7x28_mod_9982(clk,rst,matrix_A[9982],matrix_B[182],mul_res1[9982]);
multi_7x28 multi_7x28_mod_9983(clk,rst,matrix_A[9983],matrix_B[183],mul_res1[9983]);
multi_7x28 multi_7x28_mod_9984(clk,rst,matrix_A[9984],matrix_B[184],mul_res1[9984]);
multi_7x28 multi_7x28_mod_9985(clk,rst,matrix_A[9985],matrix_B[185],mul_res1[9985]);
multi_7x28 multi_7x28_mod_9986(clk,rst,matrix_A[9986],matrix_B[186],mul_res1[9986]);
multi_7x28 multi_7x28_mod_9987(clk,rst,matrix_A[9987],matrix_B[187],mul_res1[9987]);
multi_7x28 multi_7x28_mod_9988(clk,rst,matrix_A[9988],matrix_B[188],mul_res1[9988]);
multi_7x28 multi_7x28_mod_9989(clk,rst,matrix_A[9989],matrix_B[189],mul_res1[9989]);
multi_7x28 multi_7x28_mod_9990(clk,rst,matrix_A[9990],matrix_B[190],mul_res1[9990]);
multi_7x28 multi_7x28_mod_9991(clk,rst,matrix_A[9991],matrix_B[191],mul_res1[9991]);
multi_7x28 multi_7x28_mod_9992(clk,rst,matrix_A[9992],matrix_B[192],mul_res1[9992]);
multi_7x28 multi_7x28_mod_9993(clk,rst,matrix_A[9993],matrix_B[193],mul_res1[9993]);
multi_7x28 multi_7x28_mod_9994(clk,rst,matrix_A[9994],matrix_B[194],mul_res1[9994]);
multi_7x28 multi_7x28_mod_9995(clk,rst,matrix_A[9995],matrix_B[195],mul_res1[9995]);
multi_7x28 multi_7x28_mod_9996(clk,rst,matrix_A[9996],matrix_B[196],mul_res1[9996]);
multi_7x28 multi_7x28_mod_9997(clk,rst,matrix_A[9997],matrix_B[197],mul_res1[9997]);
multi_7x28 multi_7x28_mod_9998(clk,rst,matrix_A[9998],matrix_B[198],mul_res1[9998]);
multi_7x28 multi_7x28_mod_9999(clk,rst,matrix_A[9999],matrix_B[199],mul_res1[9999]);
multi_7x28 multi_7x28_mod_10000(clk,rst,matrix_A[10000],matrix_B[0],mul_res1[10000]);
multi_7x28 multi_7x28_mod_10001(clk,rst,matrix_A[10001],matrix_B[1],mul_res1[10001]);
multi_7x28 multi_7x28_mod_10002(clk,rst,matrix_A[10002],matrix_B[2],mul_res1[10002]);
multi_7x28 multi_7x28_mod_10003(clk,rst,matrix_A[10003],matrix_B[3],mul_res1[10003]);
multi_7x28 multi_7x28_mod_10004(clk,rst,matrix_A[10004],matrix_B[4],mul_res1[10004]);
multi_7x28 multi_7x28_mod_10005(clk,rst,matrix_A[10005],matrix_B[5],mul_res1[10005]);
multi_7x28 multi_7x28_mod_10006(clk,rst,matrix_A[10006],matrix_B[6],mul_res1[10006]);
multi_7x28 multi_7x28_mod_10007(clk,rst,matrix_A[10007],matrix_B[7],mul_res1[10007]);
multi_7x28 multi_7x28_mod_10008(clk,rst,matrix_A[10008],matrix_B[8],mul_res1[10008]);
multi_7x28 multi_7x28_mod_10009(clk,rst,matrix_A[10009],matrix_B[9],mul_res1[10009]);
multi_7x28 multi_7x28_mod_10010(clk,rst,matrix_A[10010],matrix_B[10],mul_res1[10010]);
multi_7x28 multi_7x28_mod_10011(clk,rst,matrix_A[10011],matrix_B[11],mul_res1[10011]);
multi_7x28 multi_7x28_mod_10012(clk,rst,matrix_A[10012],matrix_B[12],mul_res1[10012]);
multi_7x28 multi_7x28_mod_10013(clk,rst,matrix_A[10013],matrix_B[13],mul_res1[10013]);
multi_7x28 multi_7x28_mod_10014(clk,rst,matrix_A[10014],matrix_B[14],mul_res1[10014]);
multi_7x28 multi_7x28_mod_10015(clk,rst,matrix_A[10015],matrix_B[15],mul_res1[10015]);
multi_7x28 multi_7x28_mod_10016(clk,rst,matrix_A[10016],matrix_B[16],mul_res1[10016]);
multi_7x28 multi_7x28_mod_10017(clk,rst,matrix_A[10017],matrix_B[17],mul_res1[10017]);
multi_7x28 multi_7x28_mod_10018(clk,rst,matrix_A[10018],matrix_B[18],mul_res1[10018]);
multi_7x28 multi_7x28_mod_10019(clk,rst,matrix_A[10019],matrix_B[19],mul_res1[10019]);
multi_7x28 multi_7x28_mod_10020(clk,rst,matrix_A[10020],matrix_B[20],mul_res1[10020]);
multi_7x28 multi_7x28_mod_10021(clk,rst,matrix_A[10021],matrix_B[21],mul_res1[10021]);
multi_7x28 multi_7x28_mod_10022(clk,rst,matrix_A[10022],matrix_B[22],mul_res1[10022]);
multi_7x28 multi_7x28_mod_10023(clk,rst,matrix_A[10023],matrix_B[23],mul_res1[10023]);
multi_7x28 multi_7x28_mod_10024(clk,rst,matrix_A[10024],matrix_B[24],mul_res1[10024]);
multi_7x28 multi_7x28_mod_10025(clk,rst,matrix_A[10025],matrix_B[25],mul_res1[10025]);
multi_7x28 multi_7x28_mod_10026(clk,rst,matrix_A[10026],matrix_B[26],mul_res1[10026]);
multi_7x28 multi_7x28_mod_10027(clk,rst,matrix_A[10027],matrix_B[27],mul_res1[10027]);
multi_7x28 multi_7x28_mod_10028(clk,rst,matrix_A[10028],matrix_B[28],mul_res1[10028]);
multi_7x28 multi_7x28_mod_10029(clk,rst,matrix_A[10029],matrix_B[29],mul_res1[10029]);
multi_7x28 multi_7x28_mod_10030(clk,rst,matrix_A[10030],matrix_B[30],mul_res1[10030]);
multi_7x28 multi_7x28_mod_10031(clk,rst,matrix_A[10031],matrix_B[31],mul_res1[10031]);
multi_7x28 multi_7x28_mod_10032(clk,rst,matrix_A[10032],matrix_B[32],mul_res1[10032]);
multi_7x28 multi_7x28_mod_10033(clk,rst,matrix_A[10033],matrix_B[33],mul_res1[10033]);
multi_7x28 multi_7x28_mod_10034(clk,rst,matrix_A[10034],matrix_B[34],mul_res1[10034]);
multi_7x28 multi_7x28_mod_10035(clk,rst,matrix_A[10035],matrix_B[35],mul_res1[10035]);
multi_7x28 multi_7x28_mod_10036(clk,rst,matrix_A[10036],matrix_B[36],mul_res1[10036]);
multi_7x28 multi_7x28_mod_10037(clk,rst,matrix_A[10037],matrix_B[37],mul_res1[10037]);
multi_7x28 multi_7x28_mod_10038(clk,rst,matrix_A[10038],matrix_B[38],mul_res1[10038]);
multi_7x28 multi_7x28_mod_10039(clk,rst,matrix_A[10039],matrix_B[39],mul_res1[10039]);
multi_7x28 multi_7x28_mod_10040(clk,rst,matrix_A[10040],matrix_B[40],mul_res1[10040]);
multi_7x28 multi_7x28_mod_10041(clk,rst,matrix_A[10041],matrix_B[41],mul_res1[10041]);
multi_7x28 multi_7x28_mod_10042(clk,rst,matrix_A[10042],matrix_B[42],mul_res1[10042]);
multi_7x28 multi_7x28_mod_10043(clk,rst,matrix_A[10043],matrix_B[43],mul_res1[10043]);
multi_7x28 multi_7x28_mod_10044(clk,rst,matrix_A[10044],matrix_B[44],mul_res1[10044]);
multi_7x28 multi_7x28_mod_10045(clk,rst,matrix_A[10045],matrix_B[45],mul_res1[10045]);
multi_7x28 multi_7x28_mod_10046(clk,rst,matrix_A[10046],matrix_B[46],mul_res1[10046]);
multi_7x28 multi_7x28_mod_10047(clk,rst,matrix_A[10047],matrix_B[47],mul_res1[10047]);
multi_7x28 multi_7x28_mod_10048(clk,rst,matrix_A[10048],matrix_B[48],mul_res1[10048]);
multi_7x28 multi_7x28_mod_10049(clk,rst,matrix_A[10049],matrix_B[49],mul_res1[10049]);
multi_7x28 multi_7x28_mod_10050(clk,rst,matrix_A[10050],matrix_B[50],mul_res1[10050]);
multi_7x28 multi_7x28_mod_10051(clk,rst,matrix_A[10051],matrix_B[51],mul_res1[10051]);
multi_7x28 multi_7x28_mod_10052(clk,rst,matrix_A[10052],matrix_B[52],mul_res1[10052]);
multi_7x28 multi_7x28_mod_10053(clk,rst,matrix_A[10053],matrix_B[53],mul_res1[10053]);
multi_7x28 multi_7x28_mod_10054(clk,rst,matrix_A[10054],matrix_B[54],mul_res1[10054]);
multi_7x28 multi_7x28_mod_10055(clk,rst,matrix_A[10055],matrix_B[55],mul_res1[10055]);
multi_7x28 multi_7x28_mod_10056(clk,rst,matrix_A[10056],matrix_B[56],mul_res1[10056]);
multi_7x28 multi_7x28_mod_10057(clk,rst,matrix_A[10057],matrix_B[57],mul_res1[10057]);
multi_7x28 multi_7x28_mod_10058(clk,rst,matrix_A[10058],matrix_B[58],mul_res1[10058]);
multi_7x28 multi_7x28_mod_10059(clk,rst,matrix_A[10059],matrix_B[59],mul_res1[10059]);
multi_7x28 multi_7x28_mod_10060(clk,rst,matrix_A[10060],matrix_B[60],mul_res1[10060]);
multi_7x28 multi_7x28_mod_10061(clk,rst,matrix_A[10061],matrix_B[61],mul_res1[10061]);
multi_7x28 multi_7x28_mod_10062(clk,rst,matrix_A[10062],matrix_B[62],mul_res1[10062]);
multi_7x28 multi_7x28_mod_10063(clk,rst,matrix_A[10063],matrix_B[63],mul_res1[10063]);
multi_7x28 multi_7x28_mod_10064(clk,rst,matrix_A[10064],matrix_B[64],mul_res1[10064]);
multi_7x28 multi_7x28_mod_10065(clk,rst,matrix_A[10065],matrix_B[65],mul_res1[10065]);
multi_7x28 multi_7x28_mod_10066(clk,rst,matrix_A[10066],matrix_B[66],mul_res1[10066]);
multi_7x28 multi_7x28_mod_10067(clk,rst,matrix_A[10067],matrix_B[67],mul_res1[10067]);
multi_7x28 multi_7x28_mod_10068(clk,rst,matrix_A[10068],matrix_B[68],mul_res1[10068]);
multi_7x28 multi_7x28_mod_10069(clk,rst,matrix_A[10069],matrix_B[69],mul_res1[10069]);
multi_7x28 multi_7x28_mod_10070(clk,rst,matrix_A[10070],matrix_B[70],mul_res1[10070]);
multi_7x28 multi_7x28_mod_10071(clk,rst,matrix_A[10071],matrix_B[71],mul_res1[10071]);
multi_7x28 multi_7x28_mod_10072(clk,rst,matrix_A[10072],matrix_B[72],mul_res1[10072]);
multi_7x28 multi_7x28_mod_10073(clk,rst,matrix_A[10073],matrix_B[73],mul_res1[10073]);
multi_7x28 multi_7x28_mod_10074(clk,rst,matrix_A[10074],matrix_B[74],mul_res1[10074]);
multi_7x28 multi_7x28_mod_10075(clk,rst,matrix_A[10075],matrix_B[75],mul_res1[10075]);
multi_7x28 multi_7x28_mod_10076(clk,rst,matrix_A[10076],matrix_B[76],mul_res1[10076]);
multi_7x28 multi_7x28_mod_10077(clk,rst,matrix_A[10077],matrix_B[77],mul_res1[10077]);
multi_7x28 multi_7x28_mod_10078(clk,rst,matrix_A[10078],matrix_B[78],mul_res1[10078]);
multi_7x28 multi_7x28_mod_10079(clk,rst,matrix_A[10079],matrix_B[79],mul_res1[10079]);
multi_7x28 multi_7x28_mod_10080(clk,rst,matrix_A[10080],matrix_B[80],mul_res1[10080]);
multi_7x28 multi_7x28_mod_10081(clk,rst,matrix_A[10081],matrix_B[81],mul_res1[10081]);
multi_7x28 multi_7x28_mod_10082(clk,rst,matrix_A[10082],matrix_B[82],mul_res1[10082]);
multi_7x28 multi_7x28_mod_10083(clk,rst,matrix_A[10083],matrix_B[83],mul_res1[10083]);
multi_7x28 multi_7x28_mod_10084(clk,rst,matrix_A[10084],matrix_B[84],mul_res1[10084]);
multi_7x28 multi_7x28_mod_10085(clk,rst,matrix_A[10085],matrix_B[85],mul_res1[10085]);
multi_7x28 multi_7x28_mod_10086(clk,rst,matrix_A[10086],matrix_B[86],mul_res1[10086]);
multi_7x28 multi_7x28_mod_10087(clk,rst,matrix_A[10087],matrix_B[87],mul_res1[10087]);
multi_7x28 multi_7x28_mod_10088(clk,rst,matrix_A[10088],matrix_B[88],mul_res1[10088]);
multi_7x28 multi_7x28_mod_10089(clk,rst,matrix_A[10089],matrix_B[89],mul_res1[10089]);
multi_7x28 multi_7x28_mod_10090(clk,rst,matrix_A[10090],matrix_B[90],mul_res1[10090]);
multi_7x28 multi_7x28_mod_10091(clk,rst,matrix_A[10091],matrix_B[91],mul_res1[10091]);
multi_7x28 multi_7x28_mod_10092(clk,rst,matrix_A[10092],matrix_B[92],mul_res1[10092]);
multi_7x28 multi_7x28_mod_10093(clk,rst,matrix_A[10093],matrix_B[93],mul_res1[10093]);
multi_7x28 multi_7x28_mod_10094(clk,rst,matrix_A[10094],matrix_B[94],mul_res1[10094]);
multi_7x28 multi_7x28_mod_10095(clk,rst,matrix_A[10095],matrix_B[95],mul_res1[10095]);
multi_7x28 multi_7x28_mod_10096(clk,rst,matrix_A[10096],matrix_B[96],mul_res1[10096]);
multi_7x28 multi_7x28_mod_10097(clk,rst,matrix_A[10097],matrix_B[97],mul_res1[10097]);
multi_7x28 multi_7x28_mod_10098(clk,rst,matrix_A[10098],matrix_B[98],mul_res1[10098]);
multi_7x28 multi_7x28_mod_10099(clk,rst,matrix_A[10099],matrix_B[99],mul_res1[10099]);
multi_7x28 multi_7x28_mod_10100(clk,rst,matrix_A[10100],matrix_B[100],mul_res1[10100]);
multi_7x28 multi_7x28_mod_10101(clk,rst,matrix_A[10101],matrix_B[101],mul_res1[10101]);
multi_7x28 multi_7x28_mod_10102(clk,rst,matrix_A[10102],matrix_B[102],mul_res1[10102]);
multi_7x28 multi_7x28_mod_10103(clk,rst,matrix_A[10103],matrix_B[103],mul_res1[10103]);
multi_7x28 multi_7x28_mod_10104(clk,rst,matrix_A[10104],matrix_B[104],mul_res1[10104]);
multi_7x28 multi_7x28_mod_10105(clk,rst,matrix_A[10105],matrix_B[105],mul_res1[10105]);
multi_7x28 multi_7x28_mod_10106(clk,rst,matrix_A[10106],matrix_B[106],mul_res1[10106]);
multi_7x28 multi_7x28_mod_10107(clk,rst,matrix_A[10107],matrix_B[107],mul_res1[10107]);
multi_7x28 multi_7x28_mod_10108(clk,rst,matrix_A[10108],matrix_B[108],mul_res1[10108]);
multi_7x28 multi_7x28_mod_10109(clk,rst,matrix_A[10109],matrix_B[109],mul_res1[10109]);
multi_7x28 multi_7x28_mod_10110(clk,rst,matrix_A[10110],matrix_B[110],mul_res1[10110]);
multi_7x28 multi_7x28_mod_10111(clk,rst,matrix_A[10111],matrix_B[111],mul_res1[10111]);
multi_7x28 multi_7x28_mod_10112(clk,rst,matrix_A[10112],matrix_B[112],mul_res1[10112]);
multi_7x28 multi_7x28_mod_10113(clk,rst,matrix_A[10113],matrix_B[113],mul_res1[10113]);
multi_7x28 multi_7x28_mod_10114(clk,rst,matrix_A[10114],matrix_B[114],mul_res1[10114]);
multi_7x28 multi_7x28_mod_10115(clk,rst,matrix_A[10115],matrix_B[115],mul_res1[10115]);
multi_7x28 multi_7x28_mod_10116(clk,rst,matrix_A[10116],matrix_B[116],mul_res1[10116]);
multi_7x28 multi_7x28_mod_10117(clk,rst,matrix_A[10117],matrix_B[117],mul_res1[10117]);
multi_7x28 multi_7x28_mod_10118(clk,rst,matrix_A[10118],matrix_B[118],mul_res1[10118]);
multi_7x28 multi_7x28_mod_10119(clk,rst,matrix_A[10119],matrix_B[119],mul_res1[10119]);
multi_7x28 multi_7x28_mod_10120(clk,rst,matrix_A[10120],matrix_B[120],mul_res1[10120]);
multi_7x28 multi_7x28_mod_10121(clk,rst,matrix_A[10121],matrix_B[121],mul_res1[10121]);
multi_7x28 multi_7x28_mod_10122(clk,rst,matrix_A[10122],matrix_B[122],mul_res1[10122]);
multi_7x28 multi_7x28_mod_10123(clk,rst,matrix_A[10123],matrix_B[123],mul_res1[10123]);
multi_7x28 multi_7x28_mod_10124(clk,rst,matrix_A[10124],matrix_B[124],mul_res1[10124]);
multi_7x28 multi_7x28_mod_10125(clk,rst,matrix_A[10125],matrix_B[125],mul_res1[10125]);
multi_7x28 multi_7x28_mod_10126(clk,rst,matrix_A[10126],matrix_B[126],mul_res1[10126]);
multi_7x28 multi_7x28_mod_10127(clk,rst,matrix_A[10127],matrix_B[127],mul_res1[10127]);
multi_7x28 multi_7x28_mod_10128(clk,rst,matrix_A[10128],matrix_B[128],mul_res1[10128]);
multi_7x28 multi_7x28_mod_10129(clk,rst,matrix_A[10129],matrix_B[129],mul_res1[10129]);
multi_7x28 multi_7x28_mod_10130(clk,rst,matrix_A[10130],matrix_B[130],mul_res1[10130]);
multi_7x28 multi_7x28_mod_10131(clk,rst,matrix_A[10131],matrix_B[131],mul_res1[10131]);
multi_7x28 multi_7x28_mod_10132(clk,rst,matrix_A[10132],matrix_B[132],mul_res1[10132]);
multi_7x28 multi_7x28_mod_10133(clk,rst,matrix_A[10133],matrix_B[133],mul_res1[10133]);
multi_7x28 multi_7x28_mod_10134(clk,rst,matrix_A[10134],matrix_B[134],mul_res1[10134]);
multi_7x28 multi_7x28_mod_10135(clk,rst,matrix_A[10135],matrix_B[135],mul_res1[10135]);
multi_7x28 multi_7x28_mod_10136(clk,rst,matrix_A[10136],matrix_B[136],mul_res1[10136]);
multi_7x28 multi_7x28_mod_10137(clk,rst,matrix_A[10137],matrix_B[137],mul_res1[10137]);
multi_7x28 multi_7x28_mod_10138(clk,rst,matrix_A[10138],matrix_B[138],mul_res1[10138]);
multi_7x28 multi_7x28_mod_10139(clk,rst,matrix_A[10139],matrix_B[139],mul_res1[10139]);
multi_7x28 multi_7x28_mod_10140(clk,rst,matrix_A[10140],matrix_B[140],mul_res1[10140]);
multi_7x28 multi_7x28_mod_10141(clk,rst,matrix_A[10141],matrix_B[141],mul_res1[10141]);
multi_7x28 multi_7x28_mod_10142(clk,rst,matrix_A[10142],matrix_B[142],mul_res1[10142]);
multi_7x28 multi_7x28_mod_10143(clk,rst,matrix_A[10143],matrix_B[143],mul_res1[10143]);
multi_7x28 multi_7x28_mod_10144(clk,rst,matrix_A[10144],matrix_B[144],mul_res1[10144]);
multi_7x28 multi_7x28_mod_10145(clk,rst,matrix_A[10145],matrix_B[145],mul_res1[10145]);
multi_7x28 multi_7x28_mod_10146(clk,rst,matrix_A[10146],matrix_B[146],mul_res1[10146]);
multi_7x28 multi_7x28_mod_10147(clk,rst,matrix_A[10147],matrix_B[147],mul_res1[10147]);
multi_7x28 multi_7x28_mod_10148(clk,rst,matrix_A[10148],matrix_B[148],mul_res1[10148]);
multi_7x28 multi_7x28_mod_10149(clk,rst,matrix_A[10149],matrix_B[149],mul_res1[10149]);
multi_7x28 multi_7x28_mod_10150(clk,rst,matrix_A[10150],matrix_B[150],mul_res1[10150]);
multi_7x28 multi_7x28_mod_10151(clk,rst,matrix_A[10151],matrix_B[151],mul_res1[10151]);
multi_7x28 multi_7x28_mod_10152(clk,rst,matrix_A[10152],matrix_B[152],mul_res1[10152]);
multi_7x28 multi_7x28_mod_10153(clk,rst,matrix_A[10153],matrix_B[153],mul_res1[10153]);
multi_7x28 multi_7x28_mod_10154(clk,rst,matrix_A[10154],matrix_B[154],mul_res1[10154]);
multi_7x28 multi_7x28_mod_10155(clk,rst,matrix_A[10155],matrix_B[155],mul_res1[10155]);
multi_7x28 multi_7x28_mod_10156(clk,rst,matrix_A[10156],matrix_B[156],mul_res1[10156]);
multi_7x28 multi_7x28_mod_10157(clk,rst,matrix_A[10157],matrix_B[157],mul_res1[10157]);
multi_7x28 multi_7x28_mod_10158(clk,rst,matrix_A[10158],matrix_B[158],mul_res1[10158]);
multi_7x28 multi_7x28_mod_10159(clk,rst,matrix_A[10159],matrix_B[159],mul_res1[10159]);
multi_7x28 multi_7x28_mod_10160(clk,rst,matrix_A[10160],matrix_B[160],mul_res1[10160]);
multi_7x28 multi_7x28_mod_10161(clk,rst,matrix_A[10161],matrix_B[161],mul_res1[10161]);
multi_7x28 multi_7x28_mod_10162(clk,rst,matrix_A[10162],matrix_B[162],mul_res1[10162]);
multi_7x28 multi_7x28_mod_10163(clk,rst,matrix_A[10163],matrix_B[163],mul_res1[10163]);
multi_7x28 multi_7x28_mod_10164(clk,rst,matrix_A[10164],matrix_B[164],mul_res1[10164]);
multi_7x28 multi_7x28_mod_10165(clk,rst,matrix_A[10165],matrix_B[165],mul_res1[10165]);
multi_7x28 multi_7x28_mod_10166(clk,rst,matrix_A[10166],matrix_B[166],mul_res1[10166]);
multi_7x28 multi_7x28_mod_10167(clk,rst,matrix_A[10167],matrix_B[167],mul_res1[10167]);
multi_7x28 multi_7x28_mod_10168(clk,rst,matrix_A[10168],matrix_B[168],mul_res1[10168]);
multi_7x28 multi_7x28_mod_10169(clk,rst,matrix_A[10169],matrix_B[169],mul_res1[10169]);
multi_7x28 multi_7x28_mod_10170(clk,rst,matrix_A[10170],matrix_B[170],mul_res1[10170]);
multi_7x28 multi_7x28_mod_10171(clk,rst,matrix_A[10171],matrix_B[171],mul_res1[10171]);
multi_7x28 multi_7x28_mod_10172(clk,rst,matrix_A[10172],matrix_B[172],mul_res1[10172]);
multi_7x28 multi_7x28_mod_10173(clk,rst,matrix_A[10173],matrix_B[173],mul_res1[10173]);
multi_7x28 multi_7x28_mod_10174(clk,rst,matrix_A[10174],matrix_B[174],mul_res1[10174]);
multi_7x28 multi_7x28_mod_10175(clk,rst,matrix_A[10175],matrix_B[175],mul_res1[10175]);
multi_7x28 multi_7x28_mod_10176(clk,rst,matrix_A[10176],matrix_B[176],mul_res1[10176]);
multi_7x28 multi_7x28_mod_10177(clk,rst,matrix_A[10177],matrix_B[177],mul_res1[10177]);
multi_7x28 multi_7x28_mod_10178(clk,rst,matrix_A[10178],matrix_B[178],mul_res1[10178]);
multi_7x28 multi_7x28_mod_10179(clk,rst,matrix_A[10179],matrix_B[179],mul_res1[10179]);
multi_7x28 multi_7x28_mod_10180(clk,rst,matrix_A[10180],matrix_B[180],mul_res1[10180]);
multi_7x28 multi_7x28_mod_10181(clk,rst,matrix_A[10181],matrix_B[181],mul_res1[10181]);
multi_7x28 multi_7x28_mod_10182(clk,rst,matrix_A[10182],matrix_B[182],mul_res1[10182]);
multi_7x28 multi_7x28_mod_10183(clk,rst,matrix_A[10183],matrix_B[183],mul_res1[10183]);
multi_7x28 multi_7x28_mod_10184(clk,rst,matrix_A[10184],matrix_B[184],mul_res1[10184]);
multi_7x28 multi_7x28_mod_10185(clk,rst,matrix_A[10185],matrix_B[185],mul_res1[10185]);
multi_7x28 multi_7x28_mod_10186(clk,rst,matrix_A[10186],matrix_B[186],mul_res1[10186]);
multi_7x28 multi_7x28_mod_10187(clk,rst,matrix_A[10187],matrix_B[187],mul_res1[10187]);
multi_7x28 multi_7x28_mod_10188(clk,rst,matrix_A[10188],matrix_B[188],mul_res1[10188]);
multi_7x28 multi_7x28_mod_10189(clk,rst,matrix_A[10189],matrix_B[189],mul_res1[10189]);
multi_7x28 multi_7x28_mod_10190(clk,rst,matrix_A[10190],matrix_B[190],mul_res1[10190]);
multi_7x28 multi_7x28_mod_10191(clk,rst,matrix_A[10191],matrix_B[191],mul_res1[10191]);
multi_7x28 multi_7x28_mod_10192(clk,rst,matrix_A[10192],matrix_B[192],mul_res1[10192]);
multi_7x28 multi_7x28_mod_10193(clk,rst,matrix_A[10193],matrix_B[193],mul_res1[10193]);
multi_7x28 multi_7x28_mod_10194(clk,rst,matrix_A[10194],matrix_B[194],mul_res1[10194]);
multi_7x28 multi_7x28_mod_10195(clk,rst,matrix_A[10195],matrix_B[195],mul_res1[10195]);
multi_7x28 multi_7x28_mod_10196(clk,rst,matrix_A[10196],matrix_B[196],mul_res1[10196]);
multi_7x28 multi_7x28_mod_10197(clk,rst,matrix_A[10197],matrix_B[197],mul_res1[10197]);
multi_7x28 multi_7x28_mod_10198(clk,rst,matrix_A[10198],matrix_B[198],mul_res1[10198]);
multi_7x28 multi_7x28_mod_10199(clk,rst,matrix_A[10199],matrix_B[199],mul_res1[10199]);
multi_7x28 multi_7x28_mod_10200(clk,rst,matrix_A[10200],matrix_B[0],mul_res1[10200]);
multi_7x28 multi_7x28_mod_10201(clk,rst,matrix_A[10201],matrix_B[1],mul_res1[10201]);
multi_7x28 multi_7x28_mod_10202(clk,rst,matrix_A[10202],matrix_B[2],mul_res1[10202]);
multi_7x28 multi_7x28_mod_10203(clk,rst,matrix_A[10203],matrix_B[3],mul_res1[10203]);
multi_7x28 multi_7x28_mod_10204(clk,rst,matrix_A[10204],matrix_B[4],mul_res1[10204]);
multi_7x28 multi_7x28_mod_10205(clk,rst,matrix_A[10205],matrix_B[5],mul_res1[10205]);
multi_7x28 multi_7x28_mod_10206(clk,rst,matrix_A[10206],matrix_B[6],mul_res1[10206]);
multi_7x28 multi_7x28_mod_10207(clk,rst,matrix_A[10207],matrix_B[7],mul_res1[10207]);
multi_7x28 multi_7x28_mod_10208(clk,rst,matrix_A[10208],matrix_B[8],mul_res1[10208]);
multi_7x28 multi_7x28_mod_10209(clk,rst,matrix_A[10209],matrix_B[9],mul_res1[10209]);
multi_7x28 multi_7x28_mod_10210(clk,rst,matrix_A[10210],matrix_B[10],mul_res1[10210]);
multi_7x28 multi_7x28_mod_10211(clk,rst,matrix_A[10211],matrix_B[11],mul_res1[10211]);
multi_7x28 multi_7x28_mod_10212(clk,rst,matrix_A[10212],matrix_B[12],mul_res1[10212]);
multi_7x28 multi_7x28_mod_10213(clk,rst,matrix_A[10213],matrix_B[13],mul_res1[10213]);
multi_7x28 multi_7x28_mod_10214(clk,rst,matrix_A[10214],matrix_B[14],mul_res1[10214]);
multi_7x28 multi_7x28_mod_10215(clk,rst,matrix_A[10215],matrix_B[15],mul_res1[10215]);
multi_7x28 multi_7x28_mod_10216(clk,rst,matrix_A[10216],matrix_B[16],mul_res1[10216]);
multi_7x28 multi_7x28_mod_10217(clk,rst,matrix_A[10217],matrix_B[17],mul_res1[10217]);
multi_7x28 multi_7x28_mod_10218(clk,rst,matrix_A[10218],matrix_B[18],mul_res1[10218]);
multi_7x28 multi_7x28_mod_10219(clk,rst,matrix_A[10219],matrix_B[19],mul_res1[10219]);
multi_7x28 multi_7x28_mod_10220(clk,rst,matrix_A[10220],matrix_B[20],mul_res1[10220]);
multi_7x28 multi_7x28_mod_10221(clk,rst,matrix_A[10221],matrix_B[21],mul_res1[10221]);
multi_7x28 multi_7x28_mod_10222(clk,rst,matrix_A[10222],matrix_B[22],mul_res1[10222]);
multi_7x28 multi_7x28_mod_10223(clk,rst,matrix_A[10223],matrix_B[23],mul_res1[10223]);
multi_7x28 multi_7x28_mod_10224(clk,rst,matrix_A[10224],matrix_B[24],mul_res1[10224]);
multi_7x28 multi_7x28_mod_10225(clk,rst,matrix_A[10225],matrix_B[25],mul_res1[10225]);
multi_7x28 multi_7x28_mod_10226(clk,rst,matrix_A[10226],matrix_B[26],mul_res1[10226]);
multi_7x28 multi_7x28_mod_10227(clk,rst,matrix_A[10227],matrix_B[27],mul_res1[10227]);
multi_7x28 multi_7x28_mod_10228(clk,rst,matrix_A[10228],matrix_B[28],mul_res1[10228]);
multi_7x28 multi_7x28_mod_10229(clk,rst,matrix_A[10229],matrix_B[29],mul_res1[10229]);
multi_7x28 multi_7x28_mod_10230(clk,rst,matrix_A[10230],matrix_B[30],mul_res1[10230]);
multi_7x28 multi_7x28_mod_10231(clk,rst,matrix_A[10231],matrix_B[31],mul_res1[10231]);
multi_7x28 multi_7x28_mod_10232(clk,rst,matrix_A[10232],matrix_B[32],mul_res1[10232]);
multi_7x28 multi_7x28_mod_10233(clk,rst,matrix_A[10233],matrix_B[33],mul_res1[10233]);
multi_7x28 multi_7x28_mod_10234(clk,rst,matrix_A[10234],matrix_B[34],mul_res1[10234]);
multi_7x28 multi_7x28_mod_10235(clk,rst,matrix_A[10235],matrix_B[35],mul_res1[10235]);
multi_7x28 multi_7x28_mod_10236(clk,rst,matrix_A[10236],matrix_B[36],mul_res1[10236]);
multi_7x28 multi_7x28_mod_10237(clk,rst,matrix_A[10237],matrix_B[37],mul_res1[10237]);
multi_7x28 multi_7x28_mod_10238(clk,rst,matrix_A[10238],matrix_B[38],mul_res1[10238]);
multi_7x28 multi_7x28_mod_10239(clk,rst,matrix_A[10239],matrix_B[39],mul_res1[10239]);
multi_7x28 multi_7x28_mod_10240(clk,rst,matrix_A[10240],matrix_B[40],mul_res1[10240]);
multi_7x28 multi_7x28_mod_10241(clk,rst,matrix_A[10241],matrix_B[41],mul_res1[10241]);
multi_7x28 multi_7x28_mod_10242(clk,rst,matrix_A[10242],matrix_B[42],mul_res1[10242]);
multi_7x28 multi_7x28_mod_10243(clk,rst,matrix_A[10243],matrix_B[43],mul_res1[10243]);
multi_7x28 multi_7x28_mod_10244(clk,rst,matrix_A[10244],matrix_B[44],mul_res1[10244]);
multi_7x28 multi_7x28_mod_10245(clk,rst,matrix_A[10245],matrix_B[45],mul_res1[10245]);
multi_7x28 multi_7x28_mod_10246(clk,rst,matrix_A[10246],matrix_B[46],mul_res1[10246]);
multi_7x28 multi_7x28_mod_10247(clk,rst,matrix_A[10247],matrix_B[47],mul_res1[10247]);
multi_7x28 multi_7x28_mod_10248(clk,rst,matrix_A[10248],matrix_B[48],mul_res1[10248]);
multi_7x28 multi_7x28_mod_10249(clk,rst,matrix_A[10249],matrix_B[49],mul_res1[10249]);
multi_7x28 multi_7x28_mod_10250(clk,rst,matrix_A[10250],matrix_B[50],mul_res1[10250]);
multi_7x28 multi_7x28_mod_10251(clk,rst,matrix_A[10251],matrix_B[51],mul_res1[10251]);
multi_7x28 multi_7x28_mod_10252(clk,rst,matrix_A[10252],matrix_B[52],mul_res1[10252]);
multi_7x28 multi_7x28_mod_10253(clk,rst,matrix_A[10253],matrix_B[53],mul_res1[10253]);
multi_7x28 multi_7x28_mod_10254(clk,rst,matrix_A[10254],matrix_B[54],mul_res1[10254]);
multi_7x28 multi_7x28_mod_10255(clk,rst,matrix_A[10255],matrix_B[55],mul_res1[10255]);
multi_7x28 multi_7x28_mod_10256(clk,rst,matrix_A[10256],matrix_B[56],mul_res1[10256]);
multi_7x28 multi_7x28_mod_10257(clk,rst,matrix_A[10257],matrix_B[57],mul_res1[10257]);
multi_7x28 multi_7x28_mod_10258(clk,rst,matrix_A[10258],matrix_B[58],mul_res1[10258]);
multi_7x28 multi_7x28_mod_10259(clk,rst,matrix_A[10259],matrix_B[59],mul_res1[10259]);
multi_7x28 multi_7x28_mod_10260(clk,rst,matrix_A[10260],matrix_B[60],mul_res1[10260]);
multi_7x28 multi_7x28_mod_10261(clk,rst,matrix_A[10261],matrix_B[61],mul_res1[10261]);
multi_7x28 multi_7x28_mod_10262(clk,rst,matrix_A[10262],matrix_B[62],mul_res1[10262]);
multi_7x28 multi_7x28_mod_10263(clk,rst,matrix_A[10263],matrix_B[63],mul_res1[10263]);
multi_7x28 multi_7x28_mod_10264(clk,rst,matrix_A[10264],matrix_B[64],mul_res1[10264]);
multi_7x28 multi_7x28_mod_10265(clk,rst,matrix_A[10265],matrix_B[65],mul_res1[10265]);
multi_7x28 multi_7x28_mod_10266(clk,rst,matrix_A[10266],matrix_B[66],mul_res1[10266]);
multi_7x28 multi_7x28_mod_10267(clk,rst,matrix_A[10267],matrix_B[67],mul_res1[10267]);
multi_7x28 multi_7x28_mod_10268(clk,rst,matrix_A[10268],matrix_B[68],mul_res1[10268]);
multi_7x28 multi_7x28_mod_10269(clk,rst,matrix_A[10269],matrix_B[69],mul_res1[10269]);
multi_7x28 multi_7x28_mod_10270(clk,rst,matrix_A[10270],matrix_B[70],mul_res1[10270]);
multi_7x28 multi_7x28_mod_10271(clk,rst,matrix_A[10271],matrix_B[71],mul_res1[10271]);
multi_7x28 multi_7x28_mod_10272(clk,rst,matrix_A[10272],matrix_B[72],mul_res1[10272]);
multi_7x28 multi_7x28_mod_10273(clk,rst,matrix_A[10273],matrix_B[73],mul_res1[10273]);
multi_7x28 multi_7x28_mod_10274(clk,rst,matrix_A[10274],matrix_B[74],mul_res1[10274]);
multi_7x28 multi_7x28_mod_10275(clk,rst,matrix_A[10275],matrix_B[75],mul_res1[10275]);
multi_7x28 multi_7x28_mod_10276(clk,rst,matrix_A[10276],matrix_B[76],mul_res1[10276]);
multi_7x28 multi_7x28_mod_10277(clk,rst,matrix_A[10277],matrix_B[77],mul_res1[10277]);
multi_7x28 multi_7x28_mod_10278(clk,rst,matrix_A[10278],matrix_B[78],mul_res1[10278]);
multi_7x28 multi_7x28_mod_10279(clk,rst,matrix_A[10279],matrix_B[79],mul_res1[10279]);
multi_7x28 multi_7x28_mod_10280(clk,rst,matrix_A[10280],matrix_B[80],mul_res1[10280]);
multi_7x28 multi_7x28_mod_10281(clk,rst,matrix_A[10281],matrix_B[81],mul_res1[10281]);
multi_7x28 multi_7x28_mod_10282(clk,rst,matrix_A[10282],matrix_B[82],mul_res1[10282]);
multi_7x28 multi_7x28_mod_10283(clk,rst,matrix_A[10283],matrix_B[83],mul_res1[10283]);
multi_7x28 multi_7x28_mod_10284(clk,rst,matrix_A[10284],matrix_B[84],mul_res1[10284]);
multi_7x28 multi_7x28_mod_10285(clk,rst,matrix_A[10285],matrix_B[85],mul_res1[10285]);
multi_7x28 multi_7x28_mod_10286(clk,rst,matrix_A[10286],matrix_B[86],mul_res1[10286]);
multi_7x28 multi_7x28_mod_10287(clk,rst,matrix_A[10287],matrix_B[87],mul_res1[10287]);
multi_7x28 multi_7x28_mod_10288(clk,rst,matrix_A[10288],matrix_B[88],mul_res1[10288]);
multi_7x28 multi_7x28_mod_10289(clk,rst,matrix_A[10289],matrix_B[89],mul_res1[10289]);
multi_7x28 multi_7x28_mod_10290(clk,rst,matrix_A[10290],matrix_B[90],mul_res1[10290]);
multi_7x28 multi_7x28_mod_10291(clk,rst,matrix_A[10291],matrix_B[91],mul_res1[10291]);
multi_7x28 multi_7x28_mod_10292(clk,rst,matrix_A[10292],matrix_B[92],mul_res1[10292]);
multi_7x28 multi_7x28_mod_10293(clk,rst,matrix_A[10293],matrix_B[93],mul_res1[10293]);
multi_7x28 multi_7x28_mod_10294(clk,rst,matrix_A[10294],matrix_B[94],mul_res1[10294]);
multi_7x28 multi_7x28_mod_10295(clk,rst,matrix_A[10295],matrix_B[95],mul_res1[10295]);
multi_7x28 multi_7x28_mod_10296(clk,rst,matrix_A[10296],matrix_B[96],mul_res1[10296]);
multi_7x28 multi_7x28_mod_10297(clk,rst,matrix_A[10297],matrix_B[97],mul_res1[10297]);
multi_7x28 multi_7x28_mod_10298(clk,rst,matrix_A[10298],matrix_B[98],mul_res1[10298]);
multi_7x28 multi_7x28_mod_10299(clk,rst,matrix_A[10299],matrix_B[99],mul_res1[10299]);
multi_7x28 multi_7x28_mod_10300(clk,rst,matrix_A[10300],matrix_B[100],mul_res1[10300]);
multi_7x28 multi_7x28_mod_10301(clk,rst,matrix_A[10301],matrix_B[101],mul_res1[10301]);
multi_7x28 multi_7x28_mod_10302(clk,rst,matrix_A[10302],matrix_B[102],mul_res1[10302]);
multi_7x28 multi_7x28_mod_10303(clk,rst,matrix_A[10303],matrix_B[103],mul_res1[10303]);
multi_7x28 multi_7x28_mod_10304(clk,rst,matrix_A[10304],matrix_B[104],mul_res1[10304]);
multi_7x28 multi_7x28_mod_10305(clk,rst,matrix_A[10305],matrix_B[105],mul_res1[10305]);
multi_7x28 multi_7x28_mod_10306(clk,rst,matrix_A[10306],matrix_B[106],mul_res1[10306]);
multi_7x28 multi_7x28_mod_10307(clk,rst,matrix_A[10307],matrix_B[107],mul_res1[10307]);
multi_7x28 multi_7x28_mod_10308(clk,rst,matrix_A[10308],matrix_B[108],mul_res1[10308]);
multi_7x28 multi_7x28_mod_10309(clk,rst,matrix_A[10309],matrix_B[109],mul_res1[10309]);
multi_7x28 multi_7x28_mod_10310(clk,rst,matrix_A[10310],matrix_B[110],mul_res1[10310]);
multi_7x28 multi_7x28_mod_10311(clk,rst,matrix_A[10311],matrix_B[111],mul_res1[10311]);
multi_7x28 multi_7x28_mod_10312(clk,rst,matrix_A[10312],matrix_B[112],mul_res1[10312]);
multi_7x28 multi_7x28_mod_10313(clk,rst,matrix_A[10313],matrix_B[113],mul_res1[10313]);
multi_7x28 multi_7x28_mod_10314(clk,rst,matrix_A[10314],matrix_B[114],mul_res1[10314]);
multi_7x28 multi_7x28_mod_10315(clk,rst,matrix_A[10315],matrix_B[115],mul_res1[10315]);
multi_7x28 multi_7x28_mod_10316(clk,rst,matrix_A[10316],matrix_B[116],mul_res1[10316]);
multi_7x28 multi_7x28_mod_10317(clk,rst,matrix_A[10317],matrix_B[117],mul_res1[10317]);
multi_7x28 multi_7x28_mod_10318(clk,rst,matrix_A[10318],matrix_B[118],mul_res1[10318]);
multi_7x28 multi_7x28_mod_10319(clk,rst,matrix_A[10319],matrix_B[119],mul_res1[10319]);
multi_7x28 multi_7x28_mod_10320(clk,rst,matrix_A[10320],matrix_B[120],mul_res1[10320]);
multi_7x28 multi_7x28_mod_10321(clk,rst,matrix_A[10321],matrix_B[121],mul_res1[10321]);
multi_7x28 multi_7x28_mod_10322(clk,rst,matrix_A[10322],matrix_B[122],mul_res1[10322]);
multi_7x28 multi_7x28_mod_10323(clk,rst,matrix_A[10323],matrix_B[123],mul_res1[10323]);
multi_7x28 multi_7x28_mod_10324(clk,rst,matrix_A[10324],matrix_B[124],mul_res1[10324]);
multi_7x28 multi_7x28_mod_10325(clk,rst,matrix_A[10325],matrix_B[125],mul_res1[10325]);
multi_7x28 multi_7x28_mod_10326(clk,rst,matrix_A[10326],matrix_B[126],mul_res1[10326]);
multi_7x28 multi_7x28_mod_10327(clk,rst,matrix_A[10327],matrix_B[127],mul_res1[10327]);
multi_7x28 multi_7x28_mod_10328(clk,rst,matrix_A[10328],matrix_B[128],mul_res1[10328]);
multi_7x28 multi_7x28_mod_10329(clk,rst,matrix_A[10329],matrix_B[129],mul_res1[10329]);
multi_7x28 multi_7x28_mod_10330(clk,rst,matrix_A[10330],matrix_B[130],mul_res1[10330]);
multi_7x28 multi_7x28_mod_10331(clk,rst,matrix_A[10331],matrix_B[131],mul_res1[10331]);
multi_7x28 multi_7x28_mod_10332(clk,rst,matrix_A[10332],matrix_B[132],mul_res1[10332]);
multi_7x28 multi_7x28_mod_10333(clk,rst,matrix_A[10333],matrix_B[133],mul_res1[10333]);
multi_7x28 multi_7x28_mod_10334(clk,rst,matrix_A[10334],matrix_B[134],mul_res1[10334]);
multi_7x28 multi_7x28_mod_10335(clk,rst,matrix_A[10335],matrix_B[135],mul_res1[10335]);
multi_7x28 multi_7x28_mod_10336(clk,rst,matrix_A[10336],matrix_B[136],mul_res1[10336]);
multi_7x28 multi_7x28_mod_10337(clk,rst,matrix_A[10337],matrix_B[137],mul_res1[10337]);
multi_7x28 multi_7x28_mod_10338(clk,rst,matrix_A[10338],matrix_B[138],mul_res1[10338]);
multi_7x28 multi_7x28_mod_10339(clk,rst,matrix_A[10339],matrix_B[139],mul_res1[10339]);
multi_7x28 multi_7x28_mod_10340(clk,rst,matrix_A[10340],matrix_B[140],mul_res1[10340]);
multi_7x28 multi_7x28_mod_10341(clk,rst,matrix_A[10341],matrix_B[141],mul_res1[10341]);
multi_7x28 multi_7x28_mod_10342(clk,rst,matrix_A[10342],matrix_B[142],mul_res1[10342]);
multi_7x28 multi_7x28_mod_10343(clk,rst,matrix_A[10343],matrix_B[143],mul_res1[10343]);
multi_7x28 multi_7x28_mod_10344(clk,rst,matrix_A[10344],matrix_B[144],mul_res1[10344]);
multi_7x28 multi_7x28_mod_10345(clk,rst,matrix_A[10345],matrix_B[145],mul_res1[10345]);
multi_7x28 multi_7x28_mod_10346(clk,rst,matrix_A[10346],matrix_B[146],mul_res1[10346]);
multi_7x28 multi_7x28_mod_10347(clk,rst,matrix_A[10347],matrix_B[147],mul_res1[10347]);
multi_7x28 multi_7x28_mod_10348(clk,rst,matrix_A[10348],matrix_B[148],mul_res1[10348]);
multi_7x28 multi_7x28_mod_10349(clk,rst,matrix_A[10349],matrix_B[149],mul_res1[10349]);
multi_7x28 multi_7x28_mod_10350(clk,rst,matrix_A[10350],matrix_B[150],mul_res1[10350]);
multi_7x28 multi_7x28_mod_10351(clk,rst,matrix_A[10351],matrix_B[151],mul_res1[10351]);
multi_7x28 multi_7x28_mod_10352(clk,rst,matrix_A[10352],matrix_B[152],mul_res1[10352]);
multi_7x28 multi_7x28_mod_10353(clk,rst,matrix_A[10353],matrix_B[153],mul_res1[10353]);
multi_7x28 multi_7x28_mod_10354(clk,rst,matrix_A[10354],matrix_B[154],mul_res1[10354]);
multi_7x28 multi_7x28_mod_10355(clk,rst,matrix_A[10355],matrix_B[155],mul_res1[10355]);
multi_7x28 multi_7x28_mod_10356(clk,rst,matrix_A[10356],matrix_B[156],mul_res1[10356]);
multi_7x28 multi_7x28_mod_10357(clk,rst,matrix_A[10357],matrix_B[157],mul_res1[10357]);
multi_7x28 multi_7x28_mod_10358(clk,rst,matrix_A[10358],matrix_B[158],mul_res1[10358]);
multi_7x28 multi_7x28_mod_10359(clk,rst,matrix_A[10359],matrix_B[159],mul_res1[10359]);
multi_7x28 multi_7x28_mod_10360(clk,rst,matrix_A[10360],matrix_B[160],mul_res1[10360]);
multi_7x28 multi_7x28_mod_10361(clk,rst,matrix_A[10361],matrix_B[161],mul_res1[10361]);
multi_7x28 multi_7x28_mod_10362(clk,rst,matrix_A[10362],matrix_B[162],mul_res1[10362]);
multi_7x28 multi_7x28_mod_10363(clk,rst,matrix_A[10363],matrix_B[163],mul_res1[10363]);
multi_7x28 multi_7x28_mod_10364(clk,rst,matrix_A[10364],matrix_B[164],mul_res1[10364]);
multi_7x28 multi_7x28_mod_10365(clk,rst,matrix_A[10365],matrix_B[165],mul_res1[10365]);
multi_7x28 multi_7x28_mod_10366(clk,rst,matrix_A[10366],matrix_B[166],mul_res1[10366]);
multi_7x28 multi_7x28_mod_10367(clk,rst,matrix_A[10367],matrix_B[167],mul_res1[10367]);
multi_7x28 multi_7x28_mod_10368(clk,rst,matrix_A[10368],matrix_B[168],mul_res1[10368]);
multi_7x28 multi_7x28_mod_10369(clk,rst,matrix_A[10369],matrix_B[169],mul_res1[10369]);
multi_7x28 multi_7x28_mod_10370(clk,rst,matrix_A[10370],matrix_B[170],mul_res1[10370]);
multi_7x28 multi_7x28_mod_10371(clk,rst,matrix_A[10371],matrix_B[171],mul_res1[10371]);
multi_7x28 multi_7x28_mod_10372(clk,rst,matrix_A[10372],matrix_B[172],mul_res1[10372]);
multi_7x28 multi_7x28_mod_10373(clk,rst,matrix_A[10373],matrix_B[173],mul_res1[10373]);
multi_7x28 multi_7x28_mod_10374(clk,rst,matrix_A[10374],matrix_B[174],mul_res1[10374]);
multi_7x28 multi_7x28_mod_10375(clk,rst,matrix_A[10375],matrix_B[175],mul_res1[10375]);
multi_7x28 multi_7x28_mod_10376(clk,rst,matrix_A[10376],matrix_B[176],mul_res1[10376]);
multi_7x28 multi_7x28_mod_10377(clk,rst,matrix_A[10377],matrix_B[177],mul_res1[10377]);
multi_7x28 multi_7x28_mod_10378(clk,rst,matrix_A[10378],matrix_B[178],mul_res1[10378]);
multi_7x28 multi_7x28_mod_10379(clk,rst,matrix_A[10379],matrix_B[179],mul_res1[10379]);
multi_7x28 multi_7x28_mod_10380(clk,rst,matrix_A[10380],matrix_B[180],mul_res1[10380]);
multi_7x28 multi_7x28_mod_10381(clk,rst,matrix_A[10381],matrix_B[181],mul_res1[10381]);
multi_7x28 multi_7x28_mod_10382(clk,rst,matrix_A[10382],matrix_B[182],mul_res1[10382]);
multi_7x28 multi_7x28_mod_10383(clk,rst,matrix_A[10383],matrix_B[183],mul_res1[10383]);
multi_7x28 multi_7x28_mod_10384(clk,rst,matrix_A[10384],matrix_B[184],mul_res1[10384]);
multi_7x28 multi_7x28_mod_10385(clk,rst,matrix_A[10385],matrix_B[185],mul_res1[10385]);
multi_7x28 multi_7x28_mod_10386(clk,rst,matrix_A[10386],matrix_B[186],mul_res1[10386]);
multi_7x28 multi_7x28_mod_10387(clk,rst,matrix_A[10387],matrix_B[187],mul_res1[10387]);
multi_7x28 multi_7x28_mod_10388(clk,rst,matrix_A[10388],matrix_B[188],mul_res1[10388]);
multi_7x28 multi_7x28_mod_10389(clk,rst,matrix_A[10389],matrix_B[189],mul_res1[10389]);
multi_7x28 multi_7x28_mod_10390(clk,rst,matrix_A[10390],matrix_B[190],mul_res1[10390]);
multi_7x28 multi_7x28_mod_10391(clk,rst,matrix_A[10391],matrix_B[191],mul_res1[10391]);
multi_7x28 multi_7x28_mod_10392(clk,rst,matrix_A[10392],matrix_B[192],mul_res1[10392]);
multi_7x28 multi_7x28_mod_10393(clk,rst,matrix_A[10393],matrix_B[193],mul_res1[10393]);
multi_7x28 multi_7x28_mod_10394(clk,rst,matrix_A[10394],matrix_B[194],mul_res1[10394]);
multi_7x28 multi_7x28_mod_10395(clk,rst,matrix_A[10395],matrix_B[195],mul_res1[10395]);
multi_7x28 multi_7x28_mod_10396(clk,rst,matrix_A[10396],matrix_B[196],mul_res1[10396]);
multi_7x28 multi_7x28_mod_10397(clk,rst,matrix_A[10397],matrix_B[197],mul_res1[10397]);
multi_7x28 multi_7x28_mod_10398(clk,rst,matrix_A[10398],matrix_B[198],mul_res1[10398]);
multi_7x28 multi_7x28_mod_10399(clk,rst,matrix_A[10399],matrix_B[199],mul_res1[10399]);
multi_7x28 multi_7x28_mod_10400(clk,rst,matrix_A[10400],matrix_B[0],mul_res1[10400]);
multi_7x28 multi_7x28_mod_10401(clk,rst,matrix_A[10401],matrix_B[1],mul_res1[10401]);
multi_7x28 multi_7x28_mod_10402(clk,rst,matrix_A[10402],matrix_B[2],mul_res1[10402]);
multi_7x28 multi_7x28_mod_10403(clk,rst,matrix_A[10403],matrix_B[3],mul_res1[10403]);
multi_7x28 multi_7x28_mod_10404(clk,rst,matrix_A[10404],matrix_B[4],mul_res1[10404]);
multi_7x28 multi_7x28_mod_10405(clk,rst,matrix_A[10405],matrix_B[5],mul_res1[10405]);
multi_7x28 multi_7x28_mod_10406(clk,rst,matrix_A[10406],matrix_B[6],mul_res1[10406]);
multi_7x28 multi_7x28_mod_10407(clk,rst,matrix_A[10407],matrix_B[7],mul_res1[10407]);
multi_7x28 multi_7x28_mod_10408(clk,rst,matrix_A[10408],matrix_B[8],mul_res1[10408]);
multi_7x28 multi_7x28_mod_10409(clk,rst,matrix_A[10409],matrix_B[9],mul_res1[10409]);
multi_7x28 multi_7x28_mod_10410(clk,rst,matrix_A[10410],matrix_B[10],mul_res1[10410]);
multi_7x28 multi_7x28_mod_10411(clk,rst,matrix_A[10411],matrix_B[11],mul_res1[10411]);
multi_7x28 multi_7x28_mod_10412(clk,rst,matrix_A[10412],matrix_B[12],mul_res1[10412]);
multi_7x28 multi_7x28_mod_10413(clk,rst,matrix_A[10413],matrix_B[13],mul_res1[10413]);
multi_7x28 multi_7x28_mod_10414(clk,rst,matrix_A[10414],matrix_B[14],mul_res1[10414]);
multi_7x28 multi_7x28_mod_10415(clk,rst,matrix_A[10415],matrix_B[15],mul_res1[10415]);
multi_7x28 multi_7x28_mod_10416(clk,rst,matrix_A[10416],matrix_B[16],mul_res1[10416]);
multi_7x28 multi_7x28_mod_10417(clk,rst,matrix_A[10417],matrix_B[17],mul_res1[10417]);
multi_7x28 multi_7x28_mod_10418(clk,rst,matrix_A[10418],matrix_B[18],mul_res1[10418]);
multi_7x28 multi_7x28_mod_10419(clk,rst,matrix_A[10419],matrix_B[19],mul_res1[10419]);
multi_7x28 multi_7x28_mod_10420(clk,rst,matrix_A[10420],matrix_B[20],mul_res1[10420]);
multi_7x28 multi_7x28_mod_10421(clk,rst,matrix_A[10421],matrix_B[21],mul_res1[10421]);
multi_7x28 multi_7x28_mod_10422(clk,rst,matrix_A[10422],matrix_B[22],mul_res1[10422]);
multi_7x28 multi_7x28_mod_10423(clk,rst,matrix_A[10423],matrix_B[23],mul_res1[10423]);
multi_7x28 multi_7x28_mod_10424(clk,rst,matrix_A[10424],matrix_B[24],mul_res1[10424]);
multi_7x28 multi_7x28_mod_10425(clk,rst,matrix_A[10425],matrix_B[25],mul_res1[10425]);
multi_7x28 multi_7x28_mod_10426(clk,rst,matrix_A[10426],matrix_B[26],mul_res1[10426]);
multi_7x28 multi_7x28_mod_10427(clk,rst,matrix_A[10427],matrix_B[27],mul_res1[10427]);
multi_7x28 multi_7x28_mod_10428(clk,rst,matrix_A[10428],matrix_B[28],mul_res1[10428]);
multi_7x28 multi_7x28_mod_10429(clk,rst,matrix_A[10429],matrix_B[29],mul_res1[10429]);
multi_7x28 multi_7x28_mod_10430(clk,rst,matrix_A[10430],matrix_B[30],mul_res1[10430]);
multi_7x28 multi_7x28_mod_10431(clk,rst,matrix_A[10431],matrix_B[31],mul_res1[10431]);
multi_7x28 multi_7x28_mod_10432(clk,rst,matrix_A[10432],matrix_B[32],mul_res1[10432]);
multi_7x28 multi_7x28_mod_10433(clk,rst,matrix_A[10433],matrix_B[33],mul_res1[10433]);
multi_7x28 multi_7x28_mod_10434(clk,rst,matrix_A[10434],matrix_B[34],mul_res1[10434]);
multi_7x28 multi_7x28_mod_10435(clk,rst,matrix_A[10435],matrix_B[35],mul_res1[10435]);
multi_7x28 multi_7x28_mod_10436(clk,rst,matrix_A[10436],matrix_B[36],mul_res1[10436]);
multi_7x28 multi_7x28_mod_10437(clk,rst,matrix_A[10437],matrix_B[37],mul_res1[10437]);
multi_7x28 multi_7x28_mod_10438(clk,rst,matrix_A[10438],matrix_B[38],mul_res1[10438]);
multi_7x28 multi_7x28_mod_10439(clk,rst,matrix_A[10439],matrix_B[39],mul_res1[10439]);
multi_7x28 multi_7x28_mod_10440(clk,rst,matrix_A[10440],matrix_B[40],mul_res1[10440]);
multi_7x28 multi_7x28_mod_10441(clk,rst,matrix_A[10441],matrix_B[41],mul_res1[10441]);
multi_7x28 multi_7x28_mod_10442(clk,rst,matrix_A[10442],matrix_B[42],mul_res1[10442]);
multi_7x28 multi_7x28_mod_10443(clk,rst,matrix_A[10443],matrix_B[43],mul_res1[10443]);
multi_7x28 multi_7x28_mod_10444(clk,rst,matrix_A[10444],matrix_B[44],mul_res1[10444]);
multi_7x28 multi_7x28_mod_10445(clk,rst,matrix_A[10445],matrix_B[45],mul_res1[10445]);
multi_7x28 multi_7x28_mod_10446(clk,rst,matrix_A[10446],matrix_B[46],mul_res1[10446]);
multi_7x28 multi_7x28_mod_10447(clk,rst,matrix_A[10447],matrix_B[47],mul_res1[10447]);
multi_7x28 multi_7x28_mod_10448(clk,rst,matrix_A[10448],matrix_B[48],mul_res1[10448]);
multi_7x28 multi_7x28_mod_10449(clk,rst,matrix_A[10449],matrix_B[49],mul_res1[10449]);
multi_7x28 multi_7x28_mod_10450(clk,rst,matrix_A[10450],matrix_B[50],mul_res1[10450]);
multi_7x28 multi_7x28_mod_10451(clk,rst,matrix_A[10451],matrix_B[51],mul_res1[10451]);
multi_7x28 multi_7x28_mod_10452(clk,rst,matrix_A[10452],matrix_B[52],mul_res1[10452]);
multi_7x28 multi_7x28_mod_10453(clk,rst,matrix_A[10453],matrix_B[53],mul_res1[10453]);
multi_7x28 multi_7x28_mod_10454(clk,rst,matrix_A[10454],matrix_B[54],mul_res1[10454]);
multi_7x28 multi_7x28_mod_10455(clk,rst,matrix_A[10455],matrix_B[55],mul_res1[10455]);
multi_7x28 multi_7x28_mod_10456(clk,rst,matrix_A[10456],matrix_B[56],mul_res1[10456]);
multi_7x28 multi_7x28_mod_10457(clk,rst,matrix_A[10457],matrix_B[57],mul_res1[10457]);
multi_7x28 multi_7x28_mod_10458(clk,rst,matrix_A[10458],matrix_B[58],mul_res1[10458]);
multi_7x28 multi_7x28_mod_10459(clk,rst,matrix_A[10459],matrix_B[59],mul_res1[10459]);
multi_7x28 multi_7x28_mod_10460(clk,rst,matrix_A[10460],matrix_B[60],mul_res1[10460]);
multi_7x28 multi_7x28_mod_10461(clk,rst,matrix_A[10461],matrix_B[61],mul_res1[10461]);
multi_7x28 multi_7x28_mod_10462(clk,rst,matrix_A[10462],matrix_B[62],mul_res1[10462]);
multi_7x28 multi_7x28_mod_10463(clk,rst,matrix_A[10463],matrix_B[63],mul_res1[10463]);
multi_7x28 multi_7x28_mod_10464(clk,rst,matrix_A[10464],matrix_B[64],mul_res1[10464]);
multi_7x28 multi_7x28_mod_10465(clk,rst,matrix_A[10465],matrix_B[65],mul_res1[10465]);
multi_7x28 multi_7x28_mod_10466(clk,rst,matrix_A[10466],matrix_B[66],mul_res1[10466]);
multi_7x28 multi_7x28_mod_10467(clk,rst,matrix_A[10467],matrix_B[67],mul_res1[10467]);
multi_7x28 multi_7x28_mod_10468(clk,rst,matrix_A[10468],matrix_B[68],mul_res1[10468]);
multi_7x28 multi_7x28_mod_10469(clk,rst,matrix_A[10469],matrix_B[69],mul_res1[10469]);
multi_7x28 multi_7x28_mod_10470(clk,rst,matrix_A[10470],matrix_B[70],mul_res1[10470]);
multi_7x28 multi_7x28_mod_10471(clk,rst,matrix_A[10471],matrix_B[71],mul_res1[10471]);
multi_7x28 multi_7x28_mod_10472(clk,rst,matrix_A[10472],matrix_B[72],mul_res1[10472]);
multi_7x28 multi_7x28_mod_10473(clk,rst,matrix_A[10473],matrix_B[73],mul_res1[10473]);
multi_7x28 multi_7x28_mod_10474(clk,rst,matrix_A[10474],matrix_B[74],mul_res1[10474]);
multi_7x28 multi_7x28_mod_10475(clk,rst,matrix_A[10475],matrix_B[75],mul_res1[10475]);
multi_7x28 multi_7x28_mod_10476(clk,rst,matrix_A[10476],matrix_B[76],mul_res1[10476]);
multi_7x28 multi_7x28_mod_10477(clk,rst,matrix_A[10477],matrix_B[77],mul_res1[10477]);
multi_7x28 multi_7x28_mod_10478(clk,rst,matrix_A[10478],matrix_B[78],mul_res1[10478]);
multi_7x28 multi_7x28_mod_10479(clk,rst,matrix_A[10479],matrix_B[79],mul_res1[10479]);
multi_7x28 multi_7x28_mod_10480(clk,rst,matrix_A[10480],matrix_B[80],mul_res1[10480]);
multi_7x28 multi_7x28_mod_10481(clk,rst,matrix_A[10481],matrix_B[81],mul_res1[10481]);
multi_7x28 multi_7x28_mod_10482(clk,rst,matrix_A[10482],matrix_B[82],mul_res1[10482]);
multi_7x28 multi_7x28_mod_10483(clk,rst,matrix_A[10483],matrix_B[83],mul_res1[10483]);
multi_7x28 multi_7x28_mod_10484(clk,rst,matrix_A[10484],matrix_B[84],mul_res1[10484]);
multi_7x28 multi_7x28_mod_10485(clk,rst,matrix_A[10485],matrix_B[85],mul_res1[10485]);
multi_7x28 multi_7x28_mod_10486(clk,rst,matrix_A[10486],matrix_B[86],mul_res1[10486]);
multi_7x28 multi_7x28_mod_10487(clk,rst,matrix_A[10487],matrix_B[87],mul_res1[10487]);
multi_7x28 multi_7x28_mod_10488(clk,rst,matrix_A[10488],matrix_B[88],mul_res1[10488]);
multi_7x28 multi_7x28_mod_10489(clk,rst,matrix_A[10489],matrix_B[89],mul_res1[10489]);
multi_7x28 multi_7x28_mod_10490(clk,rst,matrix_A[10490],matrix_B[90],mul_res1[10490]);
multi_7x28 multi_7x28_mod_10491(clk,rst,matrix_A[10491],matrix_B[91],mul_res1[10491]);
multi_7x28 multi_7x28_mod_10492(clk,rst,matrix_A[10492],matrix_B[92],mul_res1[10492]);
multi_7x28 multi_7x28_mod_10493(clk,rst,matrix_A[10493],matrix_B[93],mul_res1[10493]);
multi_7x28 multi_7x28_mod_10494(clk,rst,matrix_A[10494],matrix_B[94],mul_res1[10494]);
multi_7x28 multi_7x28_mod_10495(clk,rst,matrix_A[10495],matrix_B[95],mul_res1[10495]);
multi_7x28 multi_7x28_mod_10496(clk,rst,matrix_A[10496],matrix_B[96],mul_res1[10496]);
multi_7x28 multi_7x28_mod_10497(clk,rst,matrix_A[10497],matrix_B[97],mul_res1[10497]);
multi_7x28 multi_7x28_mod_10498(clk,rst,matrix_A[10498],matrix_B[98],mul_res1[10498]);
multi_7x28 multi_7x28_mod_10499(clk,rst,matrix_A[10499],matrix_B[99],mul_res1[10499]);
multi_7x28 multi_7x28_mod_10500(clk,rst,matrix_A[10500],matrix_B[100],mul_res1[10500]);
multi_7x28 multi_7x28_mod_10501(clk,rst,matrix_A[10501],matrix_B[101],mul_res1[10501]);
multi_7x28 multi_7x28_mod_10502(clk,rst,matrix_A[10502],matrix_B[102],mul_res1[10502]);
multi_7x28 multi_7x28_mod_10503(clk,rst,matrix_A[10503],matrix_B[103],mul_res1[10503]);
multi_7x28 multi_7x28_mod_10504(clk,rst,matrix_A[10504],matrix_B[104],mul_res1[10504]);
multi_7x28 multi_7x28_mod_10505(clk,rst,matrix_A[10505],matrix_B[105],mul_res1[10505]);
multi_7x28 multi_7x28_mod_10506(clk,rst,matrix_A[10506],matrix_B[106],mul_res1[10506]);
multi_7x28 multi_7x28_mod_10507(clk,rst,matrix_A[10507],matrix_B[107],mul_res1[10507]);
multi_7x28 multi_7x28_mod_10508(clk,rst,matrix_A[10508],matrix_B[108],mul_res1[10508]);
multi_7x28 multi_7x28_mod_10509(clk,rst,matrix_A[10509],matrix_B[109],mul_res1[10509]);
multi_7x28 multi_7x28_mod_10510(clk,rst,matrix_A[10510],matrix_B[110],mul_res1[10510]);
multi_7x28 multi_7x28_mod_10511(clk,rst,matrix_A[10511],matrix_B[111],mul_res1[10511]);
multi_7x28 multi_7x28_mod_10512(clk,rst,matrix_A[10512],matrix_B[112],mul_res1[10512]);
multi_7x28 multi_7x28_mod_10513(clk,rst,matrix_A[10513],matrix_B[113],mul_res1[10513]);
multi_7x28 multi_7x28_mod_10514(clk,rst,matrix_A[10514],matrix_B[114],mul_res1[10514]);
multi_7x28 multi_7x28_mod_10515(clk,rst,matrix_A[10515],matrix_B[115],mul_res1[10515]);
multi_7x28 multi_7x28_mod_10516(clk,rst,matrix_A[10516],matrix_B[116],mul_res1[10516]);
multi_7x28 multi_7x28_mod_10517(clk,rst,matrix_A[10517],matrix_B[117],mul_res1[10517]);
multi_7x28 multi_7x28_mod_10518(clk,rst,matrix_A[10518],matrix_B[118],mul_res1[10518]);
multi_7x28 multi_7x28_mod_10519(clk,rst,matrix_A[10519],matrix_B[119],mul_res1[10519]);
multi_7x28 multi_7x28_mod_10520(clk,rst,matrix_A[10520],matrix_B[120],mul_res1[10520]);
multi_7x28 multi_7x28_mod_10521(clk,rst,matrix_A[10521],matrix_B[121],mul_res1[10521]);
multi_7x28 multi_7x28_mod_10522(clk,rst,matrix_A[10522],matrix_B[122],mul_res1[10522]);
multi_7x28 multi_7x28_mod_10523(clk,rst,matrix_A[10523],matrix_B[123],mul_res1[10523]);
multi_7x28 multi_7x28_mod_10524(clk,rst,matrix_A[10524],matrix_B[124],mul_res1[10524]);
multi_7x28 multi_7x28_mod_10525(clk,rst,matrix_A[10525],matrix_B[125],mul_res1[10525]);
multi_7x28 multi_7x28_mod_10526(clk,rst,matrix_A[10526],matrix_B[126],mul_res1[10526]);
multi_7x28 multi_7x28_mod_10527(clk,rst,matrix_A[10527],matrix_B[127],mul_res1[10527]);
multi_7x28 multi_7x28_mod_10528(clk,rst,matrix_A[10528],matrix_B[128],mul_res1[10528]);
multi_7x28 multi_7x28_mod_10529(clk,rst,matrix_A[10529],matrix_B[129],mul_res1[10529]);
multi_7x28 multi_7x28_mod_10530(clk,rst,matrix_A[10530],matrix_B[130],mul_res1[10530]);
multi_7x28 multi_7x28_mod_10531(clk,rst,matrix_A[10531],matrix_B[131],mul_res1[10531]);
multi_7x28 multi_7x28_mod_10532(clk,rst,matrix_A[10532],matrix_B[132],mul_res1[10532]);
multi_7x28 multi_7x28_mod_10533(clk,rst,matrix_A[10533],matrix_B[133],mul_res1[10533]);
multi_7x28 multi_7x28_mod_10534(clk,rst,matrix_A[10534],matrix_B[134],mul_res1[10534]);
multi_7x28 multi_7x28_mod_10535(clk,rst,matrix_A[10535],matrix_B[135],mul_res1[10535]);
multi_7x28 multi_7x28_mod_10536(clk,rst,matrix_A[10536],matrix_B[136],mul_res1[10536]);
multi_7x28 multi_7x28_mod_10537(clk,rst,matrix_A[10537],matrix_B[137],mul_res1[10537]);
multi_7x28 multi_7x28_mod_10538(clk,rst,matrix_A[10538],matrix_B[138],mul_res1[10538]);
multi_7x28 multi_7x28_mod_10539(clk,rst,matrix_A[10539],matrix_B[139],mul_res1[10539]);
multi_7x28 multi_7x28_mod_10540(clk,rst,matrix_A[10540],matrix_B[140],mul_res1[10540]);
multi_7x28 multi_7x28_mod_10541(clk,rst,matrix_A[10541],matrix_B[141],mul_res1[10541]);
multi_7x28 multi_7x28_mod_10542(clk,rst,matrix_A[10542],matrix_B[142],mul_res1[10542]);
multi_7x28 multi_7x28_mod_10543(clk,rst,matrix_A[10543],matrix_B[143],mul_res1[10543]);
multi_7x28 multi_7x28_mod_10544(clk,rst,matrix_A[10544],matrix_B[144],mul_res1[10544]);
multi_7x28 multi_7x28_mod_10545(clk,rst,matrix_A[10545],matrix_B[145],mul_res1[10545]);
multi_7x28 multi_7x28_mod_10546(clk,rst,matrix_A[10546],matrix_B[146],mul_res1[10546]);
multi_7x28 multi_7x28_mod_10547(clk,rst,matrix_A[10547],matrix_B[147],mul_res1[10547]);
multi_7x28 multi_7x28_mod_10548(clk,rst,matrix_A[10548],matrix_B[148],mul_res1[10548]);
multi_7x28 multi_7x28_mod_10549(clk,rst,matrix_A[10549],matrix_B[149],mul_res1[10549]);
multi_7x28 multi_7x28_mod_10550(clk,rst,matrix_A[10550],matrix_B[150],mul_res1[10550]);
multi_7x28 multi_7x28_mod_10551(clk,rst,matrix_A[10551],matrix_B[151],mul_res1[10551]);
multi_7x28 multi_7x28_mod_10552(clk,rst,matrix_A[10552],matrix_B[152],mul_res1[10552]);
multi_7x28 multi_7x28_mod_10553(clk,rst,matrix_A[10553],matrix_B[153],mul_res1[10553]);
multi_7x28 multi_7x28_mod_10554(clk,rst,matrix_A[10554],matrix_B[154],mul_res1[10554]);
multi_7x28 multi_7x28_mod_10555(clk,rst,matrix_A[10555],matrix_B[155],mul_res1[10555]);
multi_7x28 multi_7x28_mod_10556(clk,rst,matrix_A[10556],matrix_B[156],mul_res1[10556]);
multi_7x28 multi_7x28_mod_10557(clk,rst,matrix_A[10557],matrix_B[157],mul_res1[10557]);
multi_7x28 multi_7x28_mod_10558(clk,rst,matrix_A[10558],matrix_B[158],mul_res1[10558]);
multi_7x28 multi_7x28_mod_10559(clk,rst,matrix_A[10559],matrix_B[159],mul_res1[10559]);
multi_7x28 multi_7x28_mod_10560(clk,rst,matrix_A[10560],matrix_B[160],mul_res1[10560]);
multi_7x28 multi_7x28_mod_10561(clk,rst,matrix_A[10561],matrix_B[161],mul_res1[10561]);
multi_7x28 multi_7x28_mod_10562(clk,rst,matrix_A[10562],matrix_B[162],mul_res1[10562]);
multi_7x28 multi_7x28_mod_10563(clk,rst,matrix_A[10563],matrix_B[163],mul_res1[10563]);
multi_7x28 multi_7x28_mod_10564(clk,rst,matrix_A[10564],matrix_B[164],mul_res1[10564]);
multi_7x28 multi_7x28_mod_10565(clk,rst,matrix_A[10565],matrix_B[165],mul_res1[10565]);
multi_7x28 multi_7x28_mod_10566(clk,rst,matrix_A[10566],matrix_B[166],mul_res1[10566]);
multi_7x28 multi_7x28_mod_10567(clk,rst,matrix_A[10567],matrix_B[167],mul_res1[10567]);
multi_7x28 multi_7x28_mod_10568(clk,rst,matrix_A[10568],matrix_B[168],mul_res1[10568]);
multi_7x28 multi_7x28_mod_10569(clk,rst,matrix_A[10569],matrix_B[169],mul_res1[10569]);
multi_7x28 multi_7x28_mod_10570(clk,rst,matrix_A[10570],matrix_B[170],mul_res1[10570]);
multi_7x28 multi_7x28_mod_10571(clk,rst,matrix_A[10571],matrix_B[171],mul_res1[10571]);
multi_7x28 multi_7x28_mod_10572(clk,rst,matrix_A[10572],matrix_B[172],mul_res1[10572]);
multi_7x28 multi_7x28_mod_10573(clk,rst,matrix_A[10573],matrix_B[173],mul_res1[10573]);
multi_7x28 multi_7x28_mod_10574(clk,rst,matrix_A[10574],matrix_B[174],mul_res1[10574]);
multi_7x28 multi_7x28_mod_10575(clk,rst,matrix_A[10575],matrix_B[175],mul_res1[10575]);
multi_7x28 multi_7x28_mod_10576(clk,rst,matrix_A[10576],matrix_B[176],mul_res1[10576]);
multi_7x28 multi_7x28_mod_10577(clk,rst,matrix_A[10577],matrix_B[177],mul_res1[10577]);
multi_7x28 multi_7x28_mod_10578(clk,rst,matrix_A[10578],matrix_B[178],mul_res1[10578]);
multi_7x28 multi_7x28_mod_10579(clk,rst,matrix_A[10579],matrix_B[179],mul_res1[10579]);
multi_7x28 multi_7x28_mod_10580(clk,rst,matrix_A[10580],matrix_B[180],mul_res1[10580]);
multi_7x28 multi_7x28_mod_10581(clk,rst,matrix_A[10581],matrix_B[181],mul_res1[10581]);
multi_7x28 multi_7x28_mod_10582(clk,rst,matrix_A[10582],matrix_B[182],mul_res1[10582]);
multi_7x28 multi_7x28_mod_10583(clk,rst,matrix_A[10583],matrix_B[183],mul_res1[10583]);
multi_7x28 multi_7x28_mod_10584(clk,rst,matrix_A[10584],matrix_B[184],mul_res1[10584]);
multi_7x28 multi_7x28_mod_10585(clk,rst,matrix_A[10585],matrix_B[185],mul_res1[10585]);
multi_7x28 multi_7x28_mod_10586(clk,rst,matrix_A[10586],matrix_B[186],mul_res1[10586]);
multi_7x28 multi_7x28_mod_10587(clk,rst,matrix_A[10587],matrix_B[187],mul_res1[10587]);
multi_7x28 multi_7x28_mod_10588(clk,rst,matrix_A[10588],matrix_B[188],mul_res1[10588]);
multi_7x28 multi_7x28_mod_10589(clk,rst,matrix_A[10589],matrix_B[189],mul_res1[10589]);
multi_7x28 multi_7x28_mod_10590(clk,rst,matrix_A[10590],matrix_B[190],mul_res1[10590]);
multi_7x28 multi_7x28_mod_10591(clk,rst,matrix_A[10591],matrix_B[191],mul_res1[10591]);
multi_7x28 multi_7x28_mod_10592(clk,rst,matrix_A[10592],matrix_B[192],mul_res1[10592]);
multi_7x28 multi_7x28_mod_10593(clk,rst,matrix_A[10593],matrix_B[193],mul_res1[10593]);
multi_7x28 multi_7x28_mod_10594(clk,rst,matrix_A[10594],matrix_B[194],mul_res1[10594]);
multi_7x28 multi_7x28_mod_10595(clk,rst,matrix_A[10595],matrix_B[195],mul_res1[10595]);
multi_7x28 multi_7x28_mod_10596(clk,rst,matrix_A[10596],matrix_B[196],mul_res1[10596]);
multi_7x28 multi_7x28_mod_10597(clk,rst,matrix_A[10597],matrix_B[197],mul_res1[10597]);
multi_7x28 multi_7x28_mod_10598(clk,rst,matrix_A[10598],matrix_B[198],mul_res1[10598]);
multi_7x28 multi_7x28_mod_10599(clk,rst,matrix_A[10599],matrix_B[199],mul_res1[10599]);
multi_7x28 multi_7x28_mod_10600(clk,rst,matrix_A[10600],matrix_B[0],mul_res1[10600]);
multi_7x28 multi_7x28_mod_10601(clk,rst,matrix_A[10601],matrix_B[1],mul_res1[10601]);
multi_7x28 multi_7x28_mod_10602(clk,rst,matrix_A[10602],matrix_B[2],mul_res1[10602]);
multi_7x28 multi_7x28_mod_10603(clk,rst,matrix_A[10603],matrix_B[3],mul_res1[10603]);
multi_7x28 multi_7x28_mod_10604(clk,rst,matrix_A[10604],matrix_B[4],mul_res1[10604]);
multi_7x28 multi_7x28_mod_10605(clk,rst,matrix_A[10605],matrix_B[5],mul_res1[10605]);
multi_7x28 multi_7x28_mod_10606(clk,rst,matrix_A[10606],matrix_B[6],mul_res1[10606]);
multi_7x28 multi_7x28_mod_10607(clk,rst,matrix_A[10607],matrix_B[7],mul_res1[10607]);
multi_7x28 multi_7x28_mod_10608(clk,rst,matrix_A[10608],matrix_B[8],mul_res1[10608]);
multi_7x28 multi_7x28_mod_10609(clk,rst,matrix_A[10609],matrix_B[9],mul_res1[10609]);
multi_7x28 multi_7x28_mod_10610(clk,rst,matrix_A[10610],matrix_B[10],mul_res1[10610]);
multi_7x28 multi_7x28_mod_10611(clk,rst,matrix_A[10611],matrix_B[11],mul_res1[10611]);
multi_7x28 multi_7x28_mod_10612(clk,rst,matrix_A[10612],matrix_B[12],mul_res1[10612]);
multi_7x28 multi_7x28_mod_10613(clk,rst,matrix_A[10613],matrix_B[13],mul_res1[10613]);
multi_7x28 multi_7x28_mod_10614(clk,rst,matrix_A[10614],matrix_B[14],mul_res1[10614]);
multi_7x28 multi_7x28_mod_10615(clk,rst,matrix_A[10615],matrix_B[15],mul_res1[10615]);
multi_7x28 multi_7x28_mod_10616(clk,rst,matrix_A[10616],matrix_B[16],mul_res1[10616]);
multi_7x28 multi_7x28_mod_10617(clk,rst,matrix_A[10617],matrix_B[17],mul_res1[10617]);
multi_7x28 multi_7x28_mod_10618(clk,rst,matrix_A[10618],matrix_B[18],mul_res1[10618]);
multi_7x28 multi_7x28_mod_10619(clk,rst,matrix_A[10619],matrix_B[19],mul_res1[10619]);
multi_7x28 multi_7x28_mod_10620(clk,rst,matrix_A[10620],matrix_B[20],mul_res1[10620]);
multi_7x28 multi_7x28_mod_10621(clk,rst,matrix_A[10621],matrix_B[21],mul_res1[10621]);
multi_7x28 multi_7x28_mod_10622(clk,rst,matrix_A[10622],matrix_B[22],mul_res1[10622]);
multi_7x28 multi_7x28_mod_10623(clk,rst,matrix_A[10623],matrix_B[23],mul_res1[10623]);
multi_7x28 multi_7x28_mod_10624(clk,rst,matrix_A[10624],matrix_B[24],mul_res1[10624]);
multi_7x28 multi_7x28_mod_10625(clk,rst,matrix_A[10625],matrix_B[25],mul_res1[10625]);
multi_7x28 multi_7x28_mod_10626(clk,rst,matrix_A[10626],matrix_B[26],mul_res1[10626]);
multi_7x28 multi_7x28_mod_10627(clk,rst,matrix_A[10627],matrix_B[27],mul_res1[10627]);
multi_7x28 multi_7x28_mod_10628(clk,rst,matrix_A[10628],matrix_B[28],mul_res1[10628]);
multi_7x28 multi_7x28_mod_10629(clk,rst,matrix_A[10629],matrix_B[29],mul_res1[10629]);
multi_7x28 multi_7x28_mod_10630(clk,rst,matrix_A[10630],matrix_B[30],mul_res1[10630]);
multi_7x28 multi_7x28_mod_10631(clk,rst,matrix_A[10631],matrix_B[31],mul_res1[10631]);
multi_7x28 multi_7x28_mod_10632(clk,rst,matrix_A[10632],matrix_B[32],mul_res1[10632]);
multi_7x28 multi_7x28_mod_10633(clk,rst,matrix_A[10633],matrix_B[33],mul_res1[10633]);
multi_7x28 multi_7x28_mod_10634(clk,rst,matrix_A[10634],matrix_B[34],mul_res1[10634]);
multi_7x28 multi_7x28_mod_10635(clk,rst,matrix_A[10635],matrix_B[35],mul_res1[10635]);
multi_7x28 multi_7x28_mod_10636(clk,rst,matrix_A[10636],matrix_B[36],mul_res1[10636]);
multi_7x28 multi_7x28_mod_10637(clk,rst,matrix_A[10637],matrix_B[37],mul_res1[10637]);
multi_7x28 multi_7x28_mod_10638(clk,rst,matrix_A[10638],matrix_B[38],mul_res1[10638]);
multi_7x28 multi_7x28_mod_10639(clk,rst,matrix_A[10639],matrix_B[39],mul_res1[10639]);
multi_7x28 multi_7x28_mod_10640(clk,rst,matrix_A[10640],matrix_B[40],mul_res1[10640]);
multi_7x28 multi_7x28_mod_10641(clk,rst,matrix_A[10641],matrix_B[41],mul_res1[10641]);
multi_7x28 multi_7x28_mod_10642(clk,rst,matrix_A[10642],matrix_B[42],mul_res1[10642]);
multi_7x28 multi_7x28_mod_10643(clk,rst,matrix_A[10643],matrix_B[43],mul_res1[10643]);
multi_7x28 multi_7x28_mod_10644(clk,rst,matrix_A[10644],matrix_B[44],mul_res1[10644]);
multi_7x28 multi_7x28_mod_10645(clk,rst,matrix_A[10645],matrix_B[45],mul_res1[10645]);
multi_7x28 multi_7x28_mod_10646(clk,rst,matrix_A[10646],matrix_B[46],mul_res1[10646]);
multi_7x28 multi_7x28_mod_10647(clk,rst,matrix_A[10647],matrix_B[47],mul_res1[10647]);
multi_7x28 multi_7x28_mod_10648(clk,rst,matrix_A[10648],matrix_B[48],mul_res1[10648]);
multi_7x28 multi_7x28_mod_10649(clk,rst,matrix_A[10649],matrix_B[49],mul_res1[10649]);
multi_7x28 multi_7x28_mod_10650(clk,rst,matrix_A[10650],matrix_B[50],mul_res1[10650]);
multi_7x28 multi_7x28_mod_10651(clk,rst,matrix_A[10651],matrix_B[51],mul_res1[10651]);
multi_7x28 multi_7x28_mod_10652(clk,rst,matrix_A[10652],matrix_B[52],mul_res1[10652]);
multi_7x28 multi_7x28_mod_10653(clk,rst,matrix_A[10653],matrix_B[53],mul_res1[10653]);
multi_7x28 multi_7x28_mod_10654(clk,rst,matrix_A[10654],matrix_B[54],mul_res1[10654]);
multi_7x28 multi_7x28_mod_10655(clk,rst,matrix_A[10655],matrix_B[55],mul_res1[10655]);
multi_7x28 multi_7x28_mod_10656(clk,rst,matrix_A[10656],matrix_B[56],mul_res1[10656]);
multi_7x28 multi_7x28_mod_10657(clk,rst,matrix_A[10657],matrix_B[57],mul_res1[10657]);
multi_7x28 multi_7x28_mod_10658(clk,rst,matrix_A[10658],matrix_B[58],mul_res1[10658]);
multi_7x28 multi_7x28_mod_10659(clk,rst,matrix_A[10659],matrix_B[59],mul_res1[10659]);
multi_7x28 multi_7x28_mod_10660(clk,rst,matrix_A[10660],matrix_B[60],mul_res1[10660]);
multi_7x28 multi_7x28_mod_10661(clk,rst,matrix_A[10661],matrix_B[61],mul_res1[10661]);
multi_7x28 multi_7x28_mod_10662(clk,rst,matrix_A[10662],matrix_B[62],mul_res1[10662]);
multi_7x28 multi_7x28_mod_10663(clk,rst,matrix_A[10663],matrix_B[63],mul_res1[10663]);
multi_7x28 multi_7x28_mod_10664(clk,rst,matrix_A[10664],matrix_B[64],mul_res1[10664]);
multi_7x28 multi_7x28_mod_10665(clk,rst,matrix_A[10665],matrix_B[65],mul_res1[10665]);
multi_7x28 multi_7x28_mod_10666(clk,rst,matrix_A[10666],matrix_B[66],mul_res1[10666]);
multi_7x28 multi_7x28_mod_10667(clk,rst,matrix_A[10667],matrix_B[67],mul_res1[10667]);
multi_7x28 multi_7x28_mod_10668(clk,rst,matrix_A[10668],matrix_B[68],mul_res1[10668]);
multi_7x28 multi_7x28_mod_10669(clk,rst,matrix_A[10669],matrix_B[69],mul_res1[10669]);
multi_7x28 multi_7x28_mod_10670(clk,rst,matrix_A[10670],matrix_B[70],mul_res1[10670]);
multi_7x28 multi_7x28_mod_10671(clk,rst,matrix_A[10671],matrix_B[71],mul_res1[10671]);
multi_7x28 multi_7x28_mod_10672(clk,rst,matrix_A[10672],matrix_B[72],mul_res1[10672]);
multi_7x28 multi_7x28_mod_10673(clk,rst,matrix_A[10673],matrix_B[73],mul_res1[10673]);
multi_7x28 multi_7x28_mod_10674(clk,rst,matrix_A[10674],matrix_B[74],mul_res1[10674]);
multi_7x28 multi_7x28_mod_10675(clk,rst,matrix_A[10675],matrix_B[75],mul_res1[10675]);
multi_7x28 multi_7x28_mod_10676(clk,rst,matrix_A[10676],matrix_B[76],mul_res1[10676]);
multi_7x28 multi_7x28_mod_10677(clk,rst,matrix_A[10677],matrix_B[77],mul_res1[10677]);
multi_7x28 multi_7x28_mod_10678(clk,rst,matrix_A[10678],matrix_B[78],mul_res1[10678]);
multi_7x28 multi_7x28_mod_10679(clk,rst,matrix_A[10679],matrix_B[79],mul_res1[10679]);
multi_7x28 multi_7x28_mod_10680(clk,rst,matrix_A[10680],matrix_B[80],mul_res1[10680]);
multi_7x28 multi_7x28_mod_10681(clk,rst,matrix_A[10681],matrix_B[81],mul_res1[10681]);
multi_7x28 multi_7x28_mod_10682(clk,rst,matrix_A[10682],matrix_B[82],mul_res1[10682]);
multi_7x28 multi_7x28_mod_10683(clk,rst,matrix_A[10683],matrix_B[83],mul_res1[10683]);
multi_7x28 multi_7x28_mod_10684(clk,rst,matrix_A[10684],matrix_B[84],mul_res1[10684]);
multi_7x28 multi_7x28_mod_10685(clk,rst,matrix_A[10685],matrix_B[85],mul_res1[10685]);
multi_7x28 multi_7x28_mod_10686(clk,rst,matrix_A[10686],matrix_B[86],mul_res1[10686]);
multi_7x28 multi_7x28_mod_10687(clk,rst,matrix_A[10687],matrix_B[87],mul_res1[10687]);
multi_7x28 multi_7x28_mod_10688(clk,rst,matrix_A[10688],matrix_B[88],mul_res1[10688]);
multi_7x28 multi_7x28_mod_10689(clk,rst,matrix_A[10689],matrix_B[89],mul_res1[10689]);
multi_7x28 multi_7x28_mod_10690(clk,rst,matrix_A[10690],matrix_B[90],mul_res1[10690]);
multi_7x28 multi_7x28_mod_10691(clk,rst,matrix_A[10691],matrix_B[91],mul_res1[10691]);
multi_7x28 multi_7x28_mod_10692(clk,rst,matrix_A[10692],matrix_B[92],mul_res1[10692]);
multi_7x28 multi_7x28_mod_10693(clk,rst,matrix_A[10693],matrix_B[93],mul_res1[10693]);
multi_7x28 multi_7x28_mod_10694(clk,rst,matrix_A[10694],matrix_B[94],mul_res1[10694]);
multi_7x28 multi_7x28_mod_10695(clk,rst,matrix_A[10695],matrix_B[95],mul_res1[10695]);
multi_7x28 multi_7x28_mod_10696(clk,rst,matrix_A[10696],matrix_B[96],mul_res1[10696]);
multi_7x28 multi_7x28_mod_10697(clk,rst,matrix_A[10697],matrix_B[97],mul_res1[10697]);
multi_7x28 multi_7x28_mod_10698(clk,rst,matrix_A[10698],matrix_B[98],mul_res1[10698]);
multi_7x28 multi_7x28_mod_10699(clk,rst,matrix_A[10699],matrix_B[99],mul_res1[10699]);
multi_7x28 multi_7x28_mod_10700(clk,rst,matrix_A[10700],matrix_B[100],mul_res1[10700]);
multi_7x28 multi_7x28_mod_10701(clk,rst,matrix_A[10701],matrix_B[101],mul_res1[10701]);
multi_7x28 multi_7x28_mod_10702(clk,rst,matrix_A[10702],matrix_B[102],mul_res1[10702]);
multi_7x28 multi_7x28_mod_10703(clk,rst,matrix_A[10703],matrix_B[103],mul_res1[10703]);
multi_7x28 multi_7x28_mod_10704(clk,rst,matrix_A[10704],matrix_B[104],mul_res1[10704]);
multi_7x28 multi_7x28_mod_10705(clk,rst,matrix_A[10705],matrix_B[105],mul_res1[10705]);
multi_7x28 multi_7x28_mod_10706(clk,rst,matrix_A[10706],matrix_B[106],mul_res1[10706]);
multi_7x28 multi_7x28_mod_10707(clk,rst,matrix_A[10707],matrix_B[107],mul_res1[10707]);
multi_7x28 multi_7x28_mod_10708(clk,rst,matrix_A[10708],matrix_B[108],mul_res1[10708]);
multi_7x28 multi_7x28_mod_10709(clk,rst,matrix_A[10709],matrix_B[109],mul_res1[10709]);
multi_7x28 multi_7x28_mod_10710(clk,rst,matrix_A[10710],matrix_B[110],mul_res1[10710]);
multi_7x28 multi_7x28_mod_10711(clk,rst,matrix_A[10711],matrix_B[111],mul_res1[10711]);
multi_7x28 multi_7x28_mod_10712(clk,rst,matrix_A[10712],matrix_B[112],mul_res1[10712]);
multi_7x28 multi_7x28_mod_10713(clk,rst,matrix_A[10713],matrix_B[113],mul_res1[10713]);
multi_7x28 multi_7x28_mod_10714(clk,rst,matrix_A[10714],matrix_B[114],mul_res1[10714]);
multi_7x28 multi_7x28_mod_10715(clk,rst,matrix_A[10715],matrix_B[115],mul_res1[10715]);
multi_7x28 multi_7x28_mod_10716(clk,rst,matrix_A[10716],matrix_B[116],mul_res1[10716]);
multi_7x28 multi_7x28_mod_10717(clk,rst,matrix_A[10717],matrix_B[117],mul_res1[10717]);
multi_7x28 multi_7x28_mod_10718(clk,rst,matrix_A[10718],matrix_B[118],mul_res1[10718]);
multi_7x28 multi_7x28_mod_10719(clk,rst,matrix_A[10719],matrix_B[119],mul_res1[10719]);
multi_7x28 multi_7x28_mod_10720(clk,rst,matrix_A[10720],matrix_B[120],mul_res1[10720]);
multi_7x28 multi_7x28_mod_10721(clk,rst,matrix_A[10721],matrix_B[121],mul_res1[10721]);
multi_7x28 multi_7x28_mod_10722(clk,rst,matrix_A[10722],matrix_B[122],mul_res1[10722]);
multi_7x28 multi_7x28_mod_10723(clk,rst,matrix_A[10723],matrix_B[123],mul_res1[10723]);
multi_7x28 multi_7x28_mod_10724(clk,rst,matrix_A[10724],matrix_B[124],mul_res1[10724]);
multi_7x28 multi_7x28_mod_10725(clk,rst,matrix_A[10725],matrix_B[125],mul_res1[10725]);
multi_7x28 multi_7x28_mod_10726(clk,rst,matrix_A[10726],matrix_B[126],mul_res1[10726]);
multi_7x28 multi_7x28_mod_10727(clk,rst,matrix_A[10727],matrix_B[127],mul_res1[10727]);
multi_7x28 multi_7x28_mod_10728(clk,rst,matrix_A[10728],matrix_B[128],mul_res1[10728]);
multi_7x28 multi_7x28_mod_10729(clk,rst,matrix_A[10729],matrix_B[129],mul_res1[10729]);
multi_7x28 multi_7x28_mod_10730(clk,rst,matrix_A[10730],matrix_B[130],mul_res1[10730]);
multi_7x28 multi_7x28_mod_10731(clk,rst,matrix_A[10731],matrix_B[131],mul_res1[10731]);
multi_7x28 multi_7x28_mod_10732(clk,rst,matrix_A[10732],matrix_B[132],mul_res1[10732]);
multi_7x28 multi_7x28_mod_10733(clk,rst,matrix_A[10733],matrix_B[133],mul_res1[10733]);
multi_7x28 multi_7x28_mod_10734(clk,rst,matrix_A[10734],matrix_B[134],mul_res1[10734]);
multi_7x28 multi_7x28_mod_10735(clk,rst,matrix_A[10735],matrix_B[135],mul_res1[10735]);
multi_7x28 multi_7x28_mod_10736(clk,rst,matrix_A[10736],matrix_B[136],mul_res1[10736]);
multi_7x28 multi_7x28_mod_10737(clk,rst,matrix_A[10737],matrix_B[137],mul_res1[10737]);
multi_7x28 multi_7x28_mod_10738(clk,rst,matrix_A[10738],matrix_B[138],mul_res1[10738]);
multi_7x28 multi_7x28_mod_10739(clk,rst,matrix_A[10739],matrix_B[139],mul_res1[10739]);
multi_7x28 multi_7x28_mod_10740(clk,rst,matrix_A[10740],matrix_B[140],mul_res1[10740]);
multi_7x28 multi_7x28_mod_10741(clk,rst,matrix_A[10741],matrix_B[141],mul_res1[10741]);
multi_7x28 multi_7x28_mod_10742(clk,rst,matrix_A[10742],matrix_B[142],mul_res1[10742]);
multi_7x28 multi_7x28_mod_10743(clk,rst,matrix_A[10743],matrix_B[143],mul_res1[10743]);
multi_7x28 multi_7x28_mod_10744(clk,rst,matrix_A[10744],matrix_B[144],mul_res1[10744]);
multi_7x28 multi_7x28_mod_10745(clk,rst,matrix_A[10745],matrix_B[145],mul_res1[10745]);
multi_7x28 multi_7x28_mod_10746(clk,rst,matrix_A[10746],matrix_B[146],mul_res1[10746]);
multi_7x28 multi_7x28_mod_10747(clk,rst,matrix_A[10747],matrix_B[147],mul_res1[10747]);
multi_7x28 multi_7x28_mod_10748(clk,rst,matrix_A[10748],matrix_B[148],mul_res1[10748]);
multi_7x28 multi_7x28_mod_10749(clk,rst,matrix_A[10749],matrix_B[149],mul_res1[10749]);
multi_7x28 multi_7x28_mod_10750(clk,rst,matrix_A[10750],matrix_B[150],mul_res1[10750]);
multi_7x28 multi_7x28_mod_10751(clk,rst,matrix_A[10751],matrix_B[151],mul_res1[10751]);
multi_7x28 multi_7x28_mod_10752(clk,rst,matrix_A[10752],matrix_B[152],mul_res1[10752]);
multi_7x28 multi_7x28_mod_10753(clk,rst,matrix_A[10753],matrix_B[153],mul_res1[10753]);
multi_7x28 multi_7x28_mod_10754(clk,rst,matrix_A[10754],matrix_B[154],mul_res1[10754]);
multi_7x28 multi_7x28_mod_10755(clk,rst,matrix_A[10755],matrix_B[155],mul_res1[10755]);
multi_7x28 multi_7x28_mod_10756(clk,rst,matrix_A[10756],matrix_B[156],mul_res1[10756]);
multi_7x28 multi_7x28_mod_10757(clk,rst,matrix_A[10757],matrix_B[157],mul_res1[10757]);
multi_7x28 multi_7x28_mod_10758(clk,rst,matrix_A[10758],matrix_B[158],mul_res1[10758]);
multi_7x28 multi_7x28_mod_10759(clk,rst,matrix_A[10759],matrix_B[159],mul_res1[10759]);
multi_7x28 multi_7x28_mod_10760(clk,rst,matrix_A[10760],matrix_B[160],mul_res1[10760]);
multi_7x28 multi_7x28_mod_10761(clk,rst,matrix_A[10761],matrix_B[161],mul_res1[10761]);
multi_7x28 multi_7x28_mod_10762(clk,rst,matrix_A[10762],matrix_B[162],mul_res1[10762]);
multi_7x28 multi_7x28_mod_10763(clk,rst,matrix_A[10763],matrix_B[163],mul_res1[10763]);
multi_7x28 multi_7x28_mod_10764(clk,rst,matrix_A[10764],matrix_B[164],mul_res1[10764]);
multi_7x28 multi_7x28_mod_10765(clk,rst,matrix_A[10765],matrix_B[165],mul_res1[10765]);
multi_7x28 multi_7x28_mod_10766(clk,rst,matrix_A[10766],matrix_B[166],mul_res1[10766]);
multi_7x28 multi_7x28_mod_10767(clk,rst,matrix_A[10767],matrix_B[167],mul_res1[10767]);
multi_7x28 multi_7x28_mod_10768(clk,rst,matrix_A[10768],matrix_B[168],mul_res1[10768]);
multi_7x28 multi_7x28_mod_10769(clk,rst,matrix_A[10769],matrix_B[169],mul_res1[10769]);
multi_7x28 multi_7x28_mod_10770(clk,rst,matrix_A[10770],matrix_B[170],mul_res1[10770]);
multi_7x28 multi_7x28_mod_10771(clk,rst,matrix_A[10771],matrix_B[171],mul_res1[10771]);
multi_7x28 multi_7x28_mod_10772(clk,rst,matrix_A[10772],matrix_B[172],mul_res1[10772]);
multi_7x28 multi_7x28_mod_10773(clk,rst,matrix_A[10773],matrix_B[173],mul_res1[10773]);
multi_7x28 multi_7x28_mod_10774(clk,rst,matrix_A[10774],matrix_B[174],mul_res1[10774]);
multi_7x28 multi_7x28_mod_10775(clk,rst,matrix_A[10775],matrix_B[175],mul_res1[10775]);
multi_7x28 multi_7x28_mod_10776(clk,rst,matrix_A[10776],matrix_B[176],mul_res1[10776]);
multi_7x28 multi_7x28_mod_10777(clk,rst,matrix_A[10777],matrix_B[177],mul_res1[10777]);
multi_7x28 multi_7x28_mod_10778(clk,rst,matrix_A[10778],matrix_B[178],mul_res1[10778]);
multi_7x28 multi_7x28_mod_10779(clk,rst,matrix_A[10779],matrix_B[179],mul_res1[10779]);
multi_7x28 multi_7x28_mod_10780(clk,rst,matrix_A[10780],matrix_B[180],mul_res1[10780]);
multi_7x28 multi_7x28_mod_10781(clk,rst,matrix_A[10781],matrix_B[181],mul_res1[10781]);
multi_7x28 multi_7x28_mod_10782(clk,rst,matrix_A[10782],matrix_B[182],mul_res1[10782]);
multi_7x28 multi_7x28_mod_10783(clk,rst,matrix_A[10783],matrix_B[183],mul_res1[10783]);
multi_7x28 multi_7x28_mod_10784(clk,rst,matrix_A[10784],matrix_B[184],mul_res1[10784]);
multi_7x28 multi_7x28_mod_10785(clk,rst,matrix_A[10785],matrix_B[185],mul_res1[10785]);
multi_7x28 multi_7x28_mod_10786(clk,rst,matrix_A[10786],matrix_B[186],mul_res1[10786]);
multi_7x28 multi_7x28_mod_10787(clk,rst,matrix_A[10787],matrix_B[187],mul_res1[10787]);
multi_7x28 multi_7x28_mod_10788(clk,rst,matrix_A[10788],matrix_B[188],mul_res1[10788]);
multi_7x28 multi_7x28_mod_10789(clk,rst,matrix_A[10789],matrix_B[189],mul_res1[10789]);
multi_7x28 multi_7x28_mod_10790(clk,rst,matrix_A[10790],matrix_B[190],mul_res1[10790]);
multi_7x28 multi_7x28_mod_10791(clk,rst,matrix_A[10791],matrix_B[191],mul_res1[10791]);
multi_7x28 multi_7x28_mod_10792(clk,rst,matrix_A[10792],matrix_B[192],mul_res1[10792]);
multi_7x28 multi_7x28_mod_10793(clk,rst,matrix_A[10793],matrix_B[193],mul_res1[10793]);
multi_7x28 multi_7x28_mod_10794(clk,rst,matrix_A[10794],matrix_B[194],mul_res1[10794]);
multi_7x28 multi_7x28_mod_10795(clk,rst,matrix_A[10795],matrix_B[195],mul_res1[10795]);
multi_7x28 multi_7x28_mod_10796(clk,rst,matrix_A[10796],matrix_B[196],mul_res1[10796]);
multi_7x28 multi_7x28_mod_10797(clk,rst,matrix_A[10797],matrix_B[197],mul_res1[10797]);
multi_7x28 multi_7x28_mod_10798(clk,rst,matrix_A[10798],matrix_B[198],mul_res1[10798]);
multi_7x28 multi_7x28_mod_10799(clk,rst,matrix_A[10799],matrix_B[199],mul_res1[10799]);
multi_7x28 multi_7x28_mod_10800(clk,rst,matrix_A[10800],matrix_B[0],mul_res1[10800]);
multi_7x28 multi_7x28_mod_10801(clk,rst,matrix_A[10801],matrix_B[1],mul_res1[10801]);
multi_7x28 multi_7x28_mod_10802(clk,rst,matrix_A[10802],matrix_B[2],mul_res1[10802]);
multi_7x28 multi_7x28_mod_10803(clk,rst,matrix_A[10803],matrix_B[3],mul_res1[10803]);
multi_7x28 multi_7x28_mod_10804(clk,rst,matrix_A[10804],matrix_B[4],mul_res1[10804]);
multi_7x28 multi_7x28_mod_10805(clk,rst,matrix_A[10805],matrix_B[5],mul_res1[10805]);
multi_7x28 multi_7x28_mod_10806(clk,rst,matrix_A[10806],matrix_B[6],mul_res1[10806]);
multi_7x28 multi_7x28_mod_10807(clk,rst,matrix_A[10807],matrix_B[7],mul_res1[10807]);
multi_7x28 multi_7x28_mod_10808(clk,rst,matrix_A[10808],matrix_B[8],mul_res1[10808]);
multi_7x28 multi_7x28_mod_10809(clk,rst,matrix_A[10809],matrix_B[9],mul_res1[10809]);
multi_7x28 multi_7x28_mod_10810(clk,rst,matrix_A[10810],matrix_B[10],mul_res1[10810]);
multi_7x28 multi_7x28_mod_10811(clk,rst,matrix_A[10811],matrix_B[11],mul_res1[10811]);
multi_7x28 multi_7x28_mod_10812(clk,rst,matrix_A[10812],matrix_B[12],mul_res1[10812]);
multi_7x28 multi_7x28_mod_10813(clk,rst,matrix_A[10813],matrix_B[13],mul_res1[10813]);
multi_7x28 multi_7x28_mod_10814(clk,rst,matrix_A[10814],matrix_B[14],mul_res1[10814]);
multi_7x28 multi_7x28_mod_10815(clk,rst,matrix_A[10815],matrix_B[15],mul_res1[10815]);
multi_7x28 multi_7x28_mod_10816(clk,rst,matrix_A[10816],matrix_B[16],mul_res1[10816]);
multi_7x28 multi_7x28_mod_10817(clk,rst,matrix_A[10817],matrix_B[17],mul_res1[10817]);
multi_7x28 multi_7x28_mod_10818(clk,rst,matrix_A[10818],matrix_B[18],mul_res1[10818]);
multi_7x28 multi_7x28_mod_10819(clk,rst,matrix_A[10819],matrix_B[19],mul_res1[10819]);
multi_7x28 multi_7x28_mod_10820(clk,rst,matrix_A[10820],matrix_B[20],mul_res1[10820]);
multi_7x28 multi_7x28_mod_10821(clk,rst,matrix_A[10821],matrix_B[21],mul_res1[10821]);
multi_7x28 multi_7x28_mod_10822(clk,rst,matrix_A[10822],matrix_B[22],mul_res1[10822]);
multi_7x28 multi_7x28_mod_10823(clk,rst,matrix_A[10823],matrix_B[23],mul_res1[10823]);
multi_7x28 multi_7x28_mod_10824(clk,rst,matrix_A[10824],matrix_B[24],mul_res1[10824]);
multi_7x28 multi_7x28_mod_10825(clk,rst,matrix_A[10825],matrix_B[25],mul_res1[10825]);
multi_7x28 multi_7x28_mod_10826(clk,rst,matrix_A[10826],matrix_B[26],mul_res1[10826]);
multi_7x28 multi_7x28_mod_10827(clk,rst,matrix_A[10827],matrix_B[27],mul_res1[10827]);
multi_7x28 multi_7x28_mod_10828(clk,rst,matrix_A[10828],matrix_B[28],mul_res1[10828]);
multi_7x28 multi_7x28_mod_10829(clk,rst,matrix_A[10829],matrix_B[29],mul_res1[10829]);
multi_7x28 multi_7x28_mod_10830(clk,rst,matrix_A[10830],matrix_B[30],mul_res1[10830]);
multi_7x28 multi_7x28_mod_10831(clk,rst,matrix_A[10831],matrix_B[31],mul_res1[10831]);
multi_7x28 multi_7x28_mod_10832(clk,rst,matrix_A[10832],matrix_B[32],mul_res1[10832]);
multi_7x28 multi_7x28_mod_10833(clk,rst,matrix_A[10833],matrix_B[33],mul_res1[10833]);
multi_7x28 multi_7x28_mod_10834(clk,rst,matrix_A[10834],matrix_B[34],mul_res1[10834]);
multi_7x28 multi_7x28_mod_10835(clk,rst,matrix_A[10835],matrix_B[35],mul_res1[10835]);
multi_7x28 multi_7x28_mod_10836(clk,rst,matrix_A[10836],matrix_B[36],mul_res1[10836]);
multi_7x28 multi_7x28_mod_10837(clk,rst,matrix_A[10837],matrix_B[37],mul_res1[10837]);
multi_7x28 multi_7x28_mod_10838(clk,rst,matrix_A[10838],matrix_B[38],mul_res1[10838]);
multi_7x28 multi_7x28_mod_10839(clk,rst,matrix_A[10839],matrix_B[39],mul_res1[10839]);
multi_7x28 multi_7x28_mod_10840(clk,rst,matrix_A[10840],matrix_B[40],mul_res1[10840]);
multi_7x28 multi_7x28_mod_10841(clk,rst,matrix_A[10841],matrix_B[41],mul_res1[10841]);
multi_7x28 multi_7x28_mod_10842(clk,rst,matrix_A[10842],matrix_B[42],mul_res1[10842]);
multi_7x28 multi_7x28_mod_10843(clk,rst,matrix_A[10843],matrix_B[43],mul_res1[10843]);
multi_7x28 multi_7x28_mod_10844(clk,rst,matrix_A[10844],matrix_B[44],mul_res1[10844]);
multi_7x28 multi_7x28_mod_10845(clk,rst,matrix_A[10845],matrix_B[45],mul_res1[10845]);
multi_7x28 multi_7x28_mod_10846(clk,rst,matrix_A[10846],matrix_B[46],mul_res1[10846]);
multi_7x28 multi_7x28_mod_10847(clk,rst,matrix_A[10847],matrix_B[47],mul_res1[10847]);
multi_7x28 multi_7x28_mod_10848(clk,rst,matrix_A[10848],matrix_B[48],mul_res1[10848]);
multi_7x28 multi_7x28_mod_10849(clk,rst,matrix_A[10849],matrix_B[49],mul_res1[10849]);
multi_7x28 multi_7x28_mod_10850(clk,rst,matrix_A[10850],matrix_B[50],mul_res1[10850]);
multi_7x28 multi_7x28_mod_10851(clk,rst,matrix_A[10851],matrix_B[51],mul_res1[10851]);
multi_7x28 multi_7x28_mod_10852(clk,rst,matrix_A[10852],matrix_B[52],mul_res1[10852]);
multi_7x28 multi_7x28_mod_10853(clk,rst,matrix_A[10853],matrix_B[53],mul_res1[10853]);
multi_7x28 multi_7x28_mod_10854(clk,rst,matrix_A[10854],matrix_B[54],mul_res1[10854]);
multi_7x28 multi_7x28_mod_10855(clk,rst,matrix_A[10855],matrix_B[55],mul_res1[10855]);
multi_7x28 multi_7x28_mod_10856(clk,rst,matrix_A[10856],matrix_B[56],mul_res1[10856]);
multi_7x28 multi_7x28_mod_10857(clk,rst,matrix_A[10857],matrix_B[57],mul_res1[10857]);
multi_7x28 multi_7x28_mod_10858(clk,rst,matrix_A[10858],matrix_B[58],mul_res1[10858]);
multi_7x28 multi_7x28_mod_10859(clk,rst,matrix_A[10859],matrix_B[59],mul_res1[10859]);
multi_7x28 multi_7x28_mod_10860(clk,rst,matrix_A[10860],matrix_B[60],mul_res1[10860]);
multi_7x28 multi_7x28_mod_10861(clk,rst,matrix_A[10861],matrix_B[61],mul_res1[10861]);
multi_7x28 multi_7x28_mod_10862(clk,rst,matrix_A[10862],matrix_B[62],mul_res1[10862]);
multi_7x28 multi_7x28_mod_10863(clk,rst,matrix_A[10863],matrix_B[63],mul_res1[10863]);
multi_7x28 multi_7x28_mod_10864(clk,rst,matrix_A[10864],matrix_B[64],mul_res1[10864]);
multi_7x28 multi_7x28_mod_10865(clk,rst,matrix_A[10865],matrix_B[65],mul_res1[10865]);
multi_7x28 multi_7x28_mod_10866(clk,rst,matrix_A[10866],matrix_B[66],mul_res1[10866]);
multi_7x28 multi_7x28_mod_10867(clk,rst,matrix_A[10867],matrix_B[67],mul_res1[10867]);
multi_7x28 multi_7x28_mod_10868(clk,rst,matrix_A[10868],matrix_B[68],mul_res1[10868]);
multi_7x28 multi_7x28_mod_10869(clk,rst,matrix_A[10869],matrix_B[69],mul_res1[10869]);
multi_7x28 multi_7x28_mod_10870(clk,rst,matrix_A[10870],matrix_B[70],mul_res1[10870]);
multi_7x28 multi_7x28_mod_10871(clk,rst,matrix_A[10871],matrix_B[71],mul_res1[10871]);
multi_7x28 multi_7x28_mod_10872(clk,rst,matrix_A[10872],matrix_B[72],mul_res1[10872]);
multi_7x28 multi_7x28_mod_10873(clk,rst,matrix_A[10873],matrix_B[73],mul_res1[10873]);
multi_7x28 multi_7x28_mod_10874(clk,rst,matrix_A[10874],matrix_B[74],mul_res1[10874]);
multi_7x28 multi_7x28_mod_10875(clk,rst,matrix_A[10875],matrix_B[75],mul_res1[10875]);
multi_7x28 multi_7x28_mod_10876(clk,rst,matrix_A[10876],matrix_B[76],mul_res1[10876]);
multi_7x28 multi_7x28_mod_10877(clk,rst,matrix_A[10877],matrix_B[77],mul_res1[10877]);
multi_7x28 multi_7x28_mod_10878(clk,rst,matrix_A[10878],matrix_B[78],mul_res1[10878]);
multi_7x28 multi_7x28_mod_10879(clk,rst,matrix_A[10879],matrix_B[79],mul_res1[10879]);
multi_7x28 multi_7x28_mod_10880(clk,rst,matrix_A[10880],matrix_B[80],mul_res1[10880]);
multi_7x28 multi_7x28_mod_10881(clk,rst,matrix_A[10881],matrix_B[81],mul_res1[10881]);
multi_7x28 multi_7x28_mod_10882(clk,rst,matrix_A[10882],matrix_B[82],mul_res1[10882]);
multi_7x28 multi_7x28_mod_10883(clk,rst,matrix_A[10883],matrix_B[83],mul_res1[10883]);
multi_7x28 multi_7x28_mod_10884(clk,rst,matrix_A[10884],matrix_B[84],mul_res1[10884]);
multi_7x28 multi_7x28_mod_10885(clk,rst,matrix_A[10885],matrix_B[85],mul_res1[10885]);
multi_7x28 multi_7x28_mod_10886(clk,rst,matrix_A[10886],matrix_B[86],mul_res1[10886]);
multi_7x28 multi_7x28_mod_10887(clk,rst,matrix_A[10887],matrix_B[87],mul_res1[10887]);
multi_7x28 multi_7x28_mod_10888(clk,rst,matrix_A[10888],matrix_B[88],mul_res1[10888]);
multi_7x28 multi_7x28_mod_10889(clk,rst,matrix_A[10889],matrix_B[89],mul_res1[10889]);
multi_7x28 multi_7x28_mod_10890(clk,rst,matrix_A[10890],matrix_B[90],mul_res1[10890]);
multi_7x28 multi_7x28_mod_10891(clk,rst,matrix_A[10891],matrix_B[91],mul_res1[10891]);
multi_7x28 multi_7x28_mod_10892(clk,rst,matrix_A[10892],matrix_B[92],mul_res1[10892]);
multi_7x28 multi_7x28_mod_10893(clk,rst,matrix_A[10893],matrix_B[93],mul_res1[10893]);
multi_7x28 multi_7x28_mod_10894(clk,rst,matrix_A[10894],matrix_B[94],mul_res1[10894]);
multi_7x28 multi_7x28_mod_10895(clk,rst,matrix_A[10895],matrix_B[95],mul_res1[10895]);
multi_7x28 multi_7x28_mod_10896(clk,rst,matrix_A[10896],matrix_B[96],mul_res1[10896]);
multi_7x28 multi_7x28_mod_10897(clk,rst,matrix_A[10897],matrix_B[97],mul_res1[10897]);
multi_7x28 multi_7x28_mod_10898(clk,rst,matrix_A[10898],matrix_B[98],mul_res1[10898]);
multi_7x28 multi_7x28_mod_10899(clk,rst,matrix_A[10899],matrix_B[99],mul_res1[10899]);
multi_7x28 multi_7x28_mod_10900(clk,rst,matrix_A[10900],matrix_B[100],mul_res1[10900]);
multi_7x28 multi_7x28_mod_10901(clk,rst,matrix_A[10901],matrix_B[101],mul_res1[10901]);
multi_7x28 multi_7x28_mod_10902(clk,rst,matrix_A[10902],matrix_B[102],mul_res1[10902]);
multi_7x28 multi_7x28_mod_10903(clk,rst,matrix_A[10903],matrix_B[103],mul_res1[10903]);
multi_7x28 multi_7x28_mod_10904(clk,rst,matrix_A[10904],matrix_B[104],mul_res1[10904]);
multi_7x28 multi_7x28_mod_10905(clk,rst,matrix_A[10905],matrix_B[105],mul_res1[10905]);
multi_7x28 multi_7x28_mod_10906(clk,rst,matrix_A[10906],matrix_B[106],mul_res1[10906]);
multi_7x28 multi_7x28_mod_10907(clk,rst,matrix_A[10907],matrix_B[107],mul_res1[10907]);
multi_7x28 multi_7x28_mod_10908(clk,rst,matrix_A[10908],matrix_B[108],mul_res1[10908]);
multi_7x28 multi_7x28_mod_10909(clk,rst,matrix_A[10909],matrix_B[109],mul_res1[10909]);
multi_7x28 multi_7x28_mod_10910(clk,rst,matrix_A[10910],matrix_B[110],mul_res1[10910]);
multi_7x28 multi_7x28_mod_10911(clk,rst,matrix_A[10911],matrix_B[111],mul_res1[10911]);
multi_7x28 multi_7x28_mod_10912(clk,rst,matrix_A[10912],matrix_B[112],mul_res1[10912]);
multi_7x28 multi_7x28_mod_10913(clk,rst,matrix_A[10913],matrix_B[113],mul_res1[10913]);
multi_7x28 multi_7x28_mod_10914(clk,rst,matrix_A[10914],matrix_B[114],mul_res1[10914]);
multi_7x28 multi_7x28_mod_10915(clk,rst,matrix_A[10915],matrix_B[115],mul_res1[10915]);
multi_7x28 multi_7x28_mod_10916(clk,rst,matrix_A[10916],matrix_B[116],mul_res1[10916]);
multi_7x28 multi_7x28_mod_10917(clk,rst,matrix_A[10917],matrix_B[117],mul_res1[10917]);
multi_7x28 multi_7x28_mod_10918(clk,rst,matrix_A[10918],matrix_B[118],mul_res1[10918]);
multi_7x28 multi_7x28_mod_10919(clk,rst,matrix_A[10919],matrix_B[119],mul_res1[10919]);
multi_7x28 multi_7x28_mod_10920(clk,rst,matrix_A[10920],matrix_B[120],mul_res1[10920]);
multi_7x28 multi_7x28_mod_10921(clk,rst,matrix_A[10921],matrix_B[121],mul_res1[10921]);
multi_7x28 multi_7x28_mod_10922(clk,rst,matrix_A[10922],matrix_B[122],mul_res1[10922]);
multi_7x28 multi_7x28_mod_10923(clk,rst,matrix_A[10923],matrix_B[123],mul_res1[10923]);
multi_7x28 multi_7x28_mod_10924(clk,rst,matrix_A[10924],matrix_B[124],mul_res1[10924]);
multi_7x28 multi_7x28_mod_10925(clk,rst,matrix_A[10925],matrix_B[125],mul_res1[10925]);
multi_7x28 multi_7x28_mod_10926(clk,rst,matrix_A[10926],matrix_B[126],mul_res1[10926]);
multi_7x28 multi_7x28_mod_10927(clk,rst,matrix_A[10927],matrix_B[127],mul_res1[10927]);
multi_7x28 multi_7x28_mod_10928(clk,rst,matrix_A[10928],matrix_B[128],mul_res1[10928]);
multi_7x28 multi_7x28_mod_10929(clk,rst,matrix_A[10929],matrix_B[129],mul_res1[10929]);
multi_7x28 multi_7x28_mod_10930(clk,rst,matrix_A[10930],matrix_B[130],mul_res1[10930]);
multi_7x28 multi_7x28_mod_10931(clk,rst,matrix_A[10931],matrix_B[131],mul_res1[10931]);
multi_7x28 multi_7x28_mod_10932(clk,rst,matrix_A[10932],matrix_B[132],mul_res1[10932]);
multi_7x28 multi_7x28_mod_10933(clk,rst,matrix_A[10933],matrix_B[133],mul_res1[10933]);
multi_7x28 multi_7x28_mod_10934(clk,rst,matrix_A[10934],matrix_B[134],mul_res1[10934]);
multi_7x28 multi_7x28_mod_10935(clk,rst,matrix_A[10935],matrix_B[135],mul_res1[10935]);
multi_7x28 multi_7x28_mod_10936(clk,rst,matrix_A[10936],matrix_B[136],mul_res1[10936]);
multi_7x28 multi_7x28_mod_10937(clk,rst,matrix_A[10937],matrix_B[137],mul_res1[10937]);
multi_7x28 multi_7x28_mod_10938(clk,rst,matrix_A[10938],matrix_B[138],mul_res1[10938]);
multi_7x28 multi_7x28_mod_10939(clk,rst,matrix_A[10939],matrix_B[139],mul_res1[10939]);
multi_7x28 multi_7x28_mod_10940(clk,rst,matrix_A[10940],matrix_B[140],mul_res1[10940]);
multi_7x28 multi_7x28_mod_10941(clk,rst,matrix_A[10941],matrix_B[141],mul_res1[10941]);
multi_7x28 multi_7x28_mod_10942(clk,rst,matrix_A[10942],matrix_B[142],mul_res1[10942]);
multi_7x28 multi_7x28_mod_10943(clk,rst,matrix_A[10943],matrix_B[143],mul_res1[10943]);
multi_7x28 multi_7x28_mod_10944(clk,rst,matrix_A[10944],matrix_B[144],mul_res1[10944]);
multi_7x28 multi_7x28_mod_10945(clk,rst,matrix_A[10945],matrix_B[145],mul_res1[10945]);
multi_7x28 multi_7x28_mod_10946(clk,rst,matrix_A[10946],matrix_B[146],mul_res1[10946]);
multi_7x28 multi_7x28_mod_10947(clk,rst,matrix_A[10947],matrix_B[147],mul_res1[10947]);
multi_7x28 multi_7x28_mod_10948(clk,rst,matrix_A[10948],matrix_B[148],mul_res1[10948]);
multi_7x28 multi_7x28_mod_10949(clk,rst,matrix_A[10949],matrix_B[149],mul_res1[10949]);
multi_7x28 multi_7x28_mod_10950(clk,rst,matrix_A[10950],matrix_B[150],mul_res1[10950]);
multi_7x28 multi_7x28_mod_10951(clk,rst,matrix_A[10951],matrix_B[151],mul_res1[10951]);
multi_7x28 multi_7x28_mod_10952(clk,rst,matrix_A[10952],matrix_B[152],mul_res1[10952]);
multi_7x28 multi_7x28_mod_10953(clk,rst,matrix_A[10953],matrix_B[153],mul_res1[10953]);
multi_7x28 multi_7x28_mod_10954(clk,rst,matrix_A[10954],matrix_B[154],mul_res1[10954]);
multi_7x28 multi_7x28_mod_10955(clk,rst,matrix_A[10955],matrix_B[155],mul_res1[10955]);
multi_7x28 multi_7x28_mod_10956(clk,rst,matrix_A[10956],matrix_B[156],mul_res1[10956]);
multi_7x28 multi_7x28_mod_10957(clk,rst,matrix_A[10957],matrix_B[157],mul_res1[10957]);
multi_7x28 multi_7x28_mod_10958(clk,rst,matrix_A[10958],matrix_B[158],mul_res1[10958]);
multi_7x28 multi_7x28_mod_10959(clk,rst,matrix_A[10959],matrix_B[159],mul_res1[10959]);
multi_7x28 multi_7x28_mod_10960(clk,rst,matrix_A[10960],matrix_B[160],mul_res1[10960]);
multi_7x28 multi_7x28_mod_10961(clk,rst,matrix_A[10961],matrix_B[161],mul_res1[10961]);
multi_7x28 multi_7x28_mod_10962(clk,rst,matrix_A[10962],matrix_B[162],mul_res1[10962]);
multi_7x28 multi_7x28_mod_10963(clk,rst,matrix_A[10963],matrix_B[163],mul_res1[10963]);
multi_7x28 multi_7x28_mod_10964(clk,rst,matrix_A[10964],matrix_B[164],mul_res1[10964]);
multi_7x28 multi_7x28_mod_10965(clk,rst,matrix_A[10965],matrix_B[165],mul_res1[10965]);
multi_7x28 multi_7x28_mod_10966(clk,rst,matrix_A[10966],matrix_B[166],mul_res1[10966]);
multi_7x28 multi_7x28_mod_10967(clk,rst,matrix_A[10967],matrix_B[167],mul_res1[10967]);
multi_7x28 multi_7x28_mod_10968(clk,rst,matrix_A[10968],matrix_B[168],mul_res1[10968]);
multi_7x28 multi_7x28_mod_10969(clk,rst,matrix_A[10969],matrix_B[169],mul_res1[10969]);
multi_7x28 multi_7x28_mod_10970(clk,rst,matrix_A[10970],matrix_B[170],mul_res1[10970]);
multi_7x28 multi_7x28_mod_10971(clk,rst,matrix_A[10971],matrix_B[171],mul_res1[10971]);
multi_7x28 multi_7x28_mod_10972(clk,rst,matrix_A[10972],matrix_B[172],mul_res1[10972]);
multi_7x28 multi_7x28_mod_10973(clk,rst,matrix_A[10973],matrix_B[173],mul_res1[10973]);
multi_7x28 multi_7x28_mod_10974(clk,rst,matrix_A[10974],matrix_B[174],mul_res1[10974]);
multi_7x28 multi_7x28_mod_10975(clk,rst,matrix_A[10975],matrix_B[175],mul_res1[10975]);
multi_7x28 multi_7x28_mod_10976(clk,rst,matrix_A[10976],matrix_B[176],mul_res1[10976]);
multi_7x28 multi_7x28_mod_10977(clk,rst,matrix_A[10977],matrix_B[177],mul_res1[10977]);
multi_7x28 multi_7x28_mod_10978(clk,rst,matrix_A[10978],matrix_B[178],mul_res1[10978]);
multi_7x28 multi_7x28_mod_10979(clk,rst,matrix_A[10979],matrix_B[179],mul_res1[10979]);
multi_7x28 multi_7x28_mod_10980(clk,rst,matrix_A[10980],matrix_B[180],mul_res1[10980]);
multi_7x28 multi_7x28_mod_10981(clk,rst,matrix_A[10981],matrix_B[181],mul_res1[10981]);
multi_7x28 multi_7x28_mod_10982(clk,rst,matrix_A[10982],matrix_B[182],mul_res1[10982]);
multi_7x28 multi_7x28_mod_10983(clk,rst,matrix_A[10983],matrix_B[183],mul_res1[10983]);
multi_7x28 multi_7x28_mod_10984(clk,rst,matrix_A[10984],matrix_B[184],mul_res1[10984]);
multi_7x28 multi_7x28_mod_10985(clk,rst,matrix_A[10985],matrix_B[185],mul_res1[10985]);
multi_7x28 multi_7x28_mod_10986(clk,rst,matrix_A[10986],matrix_B[186],mul_res1[10986]);
multi_7x28 multi_7x28_mod_10987(clk,rst,matrix_A[10987],matrix_B[187],mul_res1[10987]);
multi_7x28 multi_7x28_mod_10988(clk,rst,matrix_A[10988],matrix_B[188],mul_res1[10988]);
multi_7x28 multi_7x28_mod_10989(clk,rst,matrix_A[10989],matrix_B[189],mul_res1[10989]);
multi_7x28 multi_7x28_mod_10990(clk,rst,matrix_A[10990],matrix_B[190],mul_res1[10990]);
multi_7x28 multi_7x28_mod_10991(clk,rst,matrix_A[10991],matrix_B[191],mul_res1[10991]);
multi_7x28 multi_7x28_mod_10992(clk,rst,matrix_A[10992],matrix_B[192],mul_res1[10992]);
multi_7x28 multi_7x28_mod_10993(clk,rst,matrix_A[10993],matrix_B[193],mul_res1[10993]);
multi_7x28 multi_7x28_mod_10994(clk,rst,matrix_A[10994],matrix_B[194],mul_res1[10994]);
multi_7x28 multi_7x28_mod_10995(clk,rst,matrix_A[10995],matrix_B[195],mul_res1[10995]);
multi_7x28 multi_7x28_mod_10996(clk,rst,matrix_A[10996],matrix_B[196],mul_res1[10996]);
multi_7x28 multi_7x28_mod_10997(clk,rst,matrix_A[10997],matrix_B[197],mul_res1[10997]);
multi_7x28 multi_7x28_mod_10998(clk,rst,matrix_A[10998],matrix_B[198],mul_res1[10998]);
multi_7x28 multi_7x28_mod_10999(clk,rst,matrix_A[10999],matrix_B[199],mul_res1[10999]);
multi_7x28 multi_7x28_mod_11000(clk,rst,matrix_A[11000],matrix_B[0],mul_res1[11000]);
multi_7x28 multi_7x28_mod_11001(clk,rst,matrix_A[11001],matrix_B[1],mul_res1[11001]);
multi_7x28 multi_7x28_mod_11002(clk,rst,matrix_A[11002],matrix_B[2],mul_res1[11002]);
multi_7x28 multi_7x28_mod_11003(clk,rst,matrix_A[11003],matrix_B[3],mul_res1[11003]);
multi_7x28 multi_7x28_mod_11004(clk,rst,matrix_A[11004],matrix_B[4],mul_res1[11004]);
multi_7x28 multi_7x28_mod_11005(clk,rst,matrix_A[11005],matrix_B[5],mul_res1[11005]);
multi_7x28 multi_7x28_mod_11006(clk,rst,matrix_A[11006],matrix_B[6],mul_res1[11006]);
multi_7x28 multi_7x28_mod_11007(clk,rst,matrix_A[11007],matrix_B[7],mul_res1[11007]);
multi_7x28 multi_7x28_mod_11008(clk,rst,matrix_A[11008],matrix_B[8],mul_res1[11008]);
multi_7x28 multi_7x28_mod_11009(clk,rst,matrix_A[11009],matrix_B[9],mul_res1[11009]);
multi_7x28 multi_7x28_mod_11010(clk,rst,matrix_A[11010],matrix_B[10],mul_res1[11010]);
multi_7x28 multi_7x28_mod_11011(clk,rst,matrix_A[11011],matrix_B[11],mul_res1[11011]);
multi_7x28 multi_7x28_mod_11012(clk,rst,matrix_A[11012],matrix_B[12],mul_res1[11012]);
multi_7x28 multi_7x28_mod_11013(clk,rst,matrix_A[11013],matrix_B[13],mul_res1[11013]);
multi_7x28 multi_7x28_mod_11014(clk,rst,matrix_A[11014],matrix_B[14],mul_res1[11014]);
multi_7x28 multi_7x28_mod_11015(clk,rst,matrix_A[11015],matrix_B[15],mul_res1[11015]);
multi_7x28 multi_7x28_mod_11016(clk,rst,matrix_A[11016],matrix_B[16],mul_res1[11016]);
multi_7x28 multi_7x28_mod_11017(clk,rst,matrix_A[11017],matrix_B[17],mul_res1[11017]);
multi_7x28 multi_7x28_mod_11018(clk,rst,matrix_A[11018],matrix_B[18],mul_res1[11018]);
multi_7x28 multi_7x28_mod_11019(clk,rst,matrix_A[11019],matrix_B[19],mul_res1[11019]);
multi_7x28 multi_7x28_mod_11020(clk,rst,matrix_A[11020],matrix_B[20],mul_res1[11020]);
multi_7x28 multi_7x28_mod_11021(clk,rst,matrix_A[11021],matrix_B[21],mul_res1[11021]);
multi_7x28 multi_7x28_mod_11022(clk,rst,matrix_A[11022],matrix_B[22],mul_res1[11022]);
multi_7x28 multi_7x28_mod_11023(clk,rst,matrix_A[11023],matrix_B[23],mul_res1[11023]);
multi_7x28 multi_7x28_mod_11024(clk,rst,matrix_A[11024],matrix_B[24],mul_res1[11024]);
multi_7x28 multi_7x28_mod_11025(clk,rst,matrix_A[11025],matrix_B[25],mul_res1[11025]);
multi_7x28 multi_7x28_mod_11026(clk,rst,matrix_A[11026],matrix_B[26],mul_res1[11026]);
multi_7x28 multi_7x28_mod_11027(clk,rst,matrix_A[11027],matrix_B[27],mul_res1[11027]);
multi_7x28 multi_7x28_mod_11028(clk,rst,matrix_A[11028],matrix_B[28],mul_res1[11028]);
multi_7x28 multi_7x28_mod_11029(clk,rst,matrix_A[11029],matrix_B[29],mul_res1[11029]);
multi_7x28 multi_7x28_mod_11030(clk,rst,matrix_A[11030],matrix_B[30],mul_res1[11030]);
multi_7x28 multi_7x28_mod_11031(clk,rst,matrix_A[11031],matrix_B[31],mul_res1[11031]);
multi_7x28 multi_7x28_mod_11032(clk,rst,matrix_A[11032],matrix_B[32],mul_res1[11032]);
multi_7x28 multi_7x28_mod_11033(clk,rst,matrix_A[11033],matrix_B[33],mul_res1[11033]);
multi_7x28 multi_7x28_mod_11034(clk,rst,matrix_A[11034],matrix_B[34],mul_res1[11034]);
multi_7x28 multi_7x28_mod_11035(clk,rst,matrix_A[11035],matrix_B[35],mul_res1[11035]);
multi_7x28 multi_7x28_mod_11036(clk,rst,matrix_A[11036],matrix_B[36],mul_res1[11036]);
multi_7x28 multi_7x28_mod_11037(clk,rst,matrix_A[11037],matrix_B[37],mul_res1[11037]);
multi_7x28 multi_7x28_mod_11038(clk,rst,matrix_A[11038],matrix_B[38],mul_res1[11038]);
multi_7x28 multi_7x28_mod_11039(clk,rst,matrix_A[11039],matrix_B[39],mul_res1[11039]);
multi_7x28 multi_7x28_mod_11040(clk,rst,matrix_A[11040],matrix_B[40],mul_res1[11040]);
multi_7x28 multi_7x28_mod_11041(clk,rst,matrix_A[11041],matrix_B[41],mul_res1[11041]);
multi_7x28 multi_7x28_mod_11042(clk,rst,matrix_A[11042],matrix_B[42],mul_res1[11042]);
multi_7x28 multi_7x28_mod_11043(clk,rst,matrix_A[11043],matrix_B[43],mul_res1[11043]);
multi_7x28 multi_7x28_mod_11044(clk,rst,matrix_A[11044],matrix_B[44],mul_res1[11044]);
multi_7x28 multi_7x28_mod_11045(clk,rst,matrix_A[11045],matrix_B[45],mul_res1[11045]);
multi_7x28 multi_7x28_mod_11046(clk,rst,matrix_A[11046],matrix_B[46],mul_res1[11046]);
multi_7x28 multi_7x28_mod_11047(clk,rst,matrix_A[11047],matrix_B[47],mul_res1[11047]);
multi_7x28 multi_7x28_mod_11048(clk,rst,matrix_A[11048],matrix_B[48],mul_res1[11048]);
multi_7x28 multi_7x28_mod_11049(clk,rst,matrix_A[11049],matrix_B[49],mul_res1[11049]);
multi_7x28 multi_7x28_mod_11050(clk,rst,matrix_A[11050],matrix_B[50],mul_res1[11050]);
multi_7x28 multi_7x28_mod_11051(clk,rst,matrix_A[11051],matrix_B[51],mul_res1[11051]);
multi_7x28 multi_7x28_mod_11052(clk,rst,matrix_A[11052],matrix_B[52],mul_res1[11052]);
multi_7x28 multi_7x28_mod_11053(clk,rst,matrix_A[11053],matrix_B[53],mul_res1[11053]);
multi_7x28 multi_7x28_mod_11054(clk,rst,matrix_A[11054],matrix_B[54],mul_res1[11054]);
multi_7x28 multi_7x28_mod_11055(clk,rst,matrix_A[11055],matrix_B[55],mul_res1[11055]);
multi_7x28 multi_7x28_mod_11056(clk,rst,matrix_A[11056],matrix_B[56],mul_res1[11056]);
multi_7x28 multi_7x28_mod_11057(clk,rst,matrix_A[11057],matrix_B[57],mul_res1[11057]);
multi_7x28 multi_7x28_mod_11058(clk,rst,matrix_A[11058],matrix_B[58],mul_res1[11058]);
multi_7x28 multi_7x28_mod_11059(clk,rst,matrix_A[11059],matrix_B[59],mul_res1[11059]);
multi_7x28 multi_7x28_mod_11060(clk,rst,matrix_A[11060],matrix_B[60],mul_res1[11060]);
multi_7x28 multi_7x28_mod_11061(clk,rst,matrix_A[11061],matrix_B[61],mul_res1[11061]);
multi_7x28 multi_7x28_mod_11062(clk,rst,matrix_A[11062],matrix_B[62],mul_res1[11062]);
multi_7x28 multi_7x28_mod_11063(clk,rst,matrix_A[11063],matrix_B[63],mul_res1[11063]);
multi_7x28 multi_7x28_mod_11064(clk,rst,matrix_A[11064],matrix_B[64],mul_res1[11064]);
multi_7x28 multi_7x28_mod_11065(clk,rst,matrix_A[11065],matrix_B[65],mul_res1[11065]);
multi_7x28 multi_7x28_mod_11066(clk,rst,matrix_A[11066],matrix_B[66],mul_res1[11066]);
multi_7x28 multi_7x28_mod_11067(clk,rst,matrix_A[11067],matrix_B[67],mul_res1[11067]);
multi_7x28 multi_7x28_mod_11068(clk,rst,matrix_A[11068],matrix_B[68],mul_res1[11068]);
multi_7x28 multi_7x28_mod_11069(clk,rst,matrix_A[11069],matrix_B[69],mul_res1[11069]);
multi_7x28 multi_7x28_mod_11070(clk,rst,matrix_A[11070],matrix_B[70],mul_res1[11070]);
multi_7x28 multi_7x28_mod_11071(clk,rst,matrix_A[11071],matrix_B[71],mul_res1[11071]);
multi_7x28 multi_7x28_mod_11072(clk,rst,matrix_A[11072],matrix_B[72],mul_res1[11072]);
multi_7x28 multi_7x28_mod_11073(clk,rst,matrix_A[11073],matrix_B[73],mul_res1[11073]);
multi_7x28 multi_7x28_mod_11074(clk,rst,matrix_A[11074],matrix_B[74],mul_res1[11074]);
multi_7x28 multi_7x28_mod_11075(clk,rst,matrix_A[11075],matrix_B[75],mul_res1[11075]);
multi_7x28 multi_7x28_mod_11076(clk,rst,matrix_A[11076],matrix_B[76],mul_res1[11076]);
multi_7x28 multi_7x28_mod_11077(clk,rst,matrix_A[11077],matrix_B[77],mul_res1[11077]);
multi_7x28 multi_7x28_mod_11078(clk,rst,matrix_A[11078],matrix_B[78],mul_res1[11078]);
multi_7x28 multi_7x28_mod_11079(clk,rst,matrix_A[11079],matrix_B[79],mul_res1[11079]);
multi_7x28 multi_7x28_mod_11080(clk,rst,matrix_A[11080],matrix_B[80],mul_res1[11080]);
multi_7x28 multi_7x28_mod_11081(clk,rst,matrix_A[11081],matrix_B[81],mul_res1[11081]);
multi_7x28 multi_7x28_mod_11082(clk,rst,matrix_A[11082],matrix_B[82],mul_res1[11082]);
multi_7x28 multi_7x28_mod_11083(clk,rst,matrix_A[11083],matrix_B[83],mul_res1[11083]);
multi_7x28 multi_7x28_mod_11084(clk,rst,matrix_A[11084],matrix_B[84],mul_res1[11084]);
multi_7x28 multi_7x28_mod_11085(clk,rst,matrix_A[11085],matrix_B[85],mul_res1[11085]);
multi_7x28 multi_7x28_mod_11086(clk,rst,matrix_A[11086],matrix_B[86],mul_res1[11086]);
multi_7x28 multi_7x28_mod_11087(clk,rst,matrix_A[11087],matrix_B[87],mul_res1[11087]);
multi_7x28 multi_7x28_mod_11088(clk,rst,matrix_A[11088],matrix_B[88],mul_res1[11088]);
multi_7x28 multi_7x28_mod_11089(clk,rst,matrix_A[11089],matrix_B[89],mul_res1[11089]);
multi_7x28 multi_7x28_mod_11090(clk,rst,matrix_A[11090],matrix_B[90],mul_res1[11090]);
multi_7x28 multi_7x28_mod_11091(clk,rst,matrix_A[11091],matrix_B[91],mul_res1[11091]);
multi_7x28 multi_7x28_mod_11092(clk,rst,matrix_A[11092],matrix_B[92],mul_res1[11092]);
multi_7x28 multi_7x28_mod_11093(clk,rst,matrix_A[11093],matrix_B[93],mul_res1[11093]);
multi_7x28 multi_7x28_mod_11094(clk,rst,matrix_A[11094],matrix_B[94],mul_res1[11094]);
multi_7x28 multi_7x28_mod_11095(clk,rst,matrix_A[11095],matrix_B[95],mul_res1[11095]);
multi_7x28 multi_7x28_mod_11096(clk,rst,matrix_A[11096],matrix_B[96],mul_res1[11096]);
multi_7x28 multi_7x28_mod_11097(clk,rst,matrix_A[11097],matrix_B[97],mul_res1[11097]);
multi_7x28 multi_7x28_mod_11098(clk,rst,matrix_A[11098],matrix_B[98],mul_res1[11098]);
multi_7x28 multi_7x28_mod_11099(clk,rst,matrix_A[11099],matrix_B[99],mul_res1[11099]);
multi_7x28 multi_7x28_mod_11100(clk,rst,matrix_A[11100],matrix_B[100],mul_res1[11100]);
multi_7x28 multi_7x28_mod_11101(clk,rst,matrix_A[11101],matrix_B[101],mul_res1[11101]);
multi_7x28 multi_7x28_mod_11102(clk,rst,matrix_A[11102],matrix_B[102],mul_res1[11102]);
multi_7x28 multi_7x28_mod_11103(clk,rst,matrix_A[11103],matrix_B[103],mul_res1[11103]);
multi_7x28 multi_7x28_mod_11104(clk,rst,matrix_A[11104],matrix_B[104],mul_res1[11104]);
multi_7x28 multi_7x28_mod_11105(clk,rst,matrix_A[11105],matrix_B[105],mul_res1[11105]);
multi_7x28 multi_7x28_mod_11106(clk,rst,matrix_A[11106],matrix_B[106],mul_res1[11106]);
multi_7x28 multi_7x28_mod_11107(clk,rst,matrix_A[11107],matrix_B[107],mul_res1[11107]);
multi_7x28 multi_7x28_mod_11108(clk,rst,matrix_A[11108],matrix_B[108],mul_res1[11108]);
multi_7x28 multi_7x28_mod_11109(clk,rst,matrix_A[11109],matrix_B[109],mul_res1[11109]);
multi_7x28 multi_7x28_mod_11110(clk,rst,matrix_A[11110],matrix_B[110],mul_res1[11110]);
multi_7x28 multi_7x28_mod_11111(clk,rst,matrix_A[11111],matrix_B[111],mul_res1[11111]);
multi_7x28 multi_7x28_mod_11112(clk,rst,matrix_A[11112],matrix_B[112],mul_res1[11112]);
multi_7x28 multi_7x28_mod_11113(clk,rst,matrix_A[11113],matrix_B[113],mul_res1[11113]);
multi_7x28 multi_7x28_mod_11114(clk,rst,matrix_A[11114],matrix_B[114],mul_res1[11114]);
multi_7x28 multi_7x28_mod_11115(clk,rst,matrix_A[11115],matrix_B[115],mul_res1[11115]);
multi_7x28 multi_7x28_mod_11116(clk,rst,matrix_A[11116],matrix_B[116],mul_res1[11116]);
multi_7x28 multi_7x28_mod_11117(clk,rst,matrix_A[11117],matrix_B[117],mul_res1[11117]);
multi_7x28 multi_7x28_mod_11118(clk,rst,matrix_A[11118],matrix_B[118],mul_res1[11118]);
multi_7x28 multi_7x28_mod_11119(clk,rst,matrix_A[11119],matrix_B[119],mul_res1[11119]);
multi_7x28 multi_7x28_mod_11120(clk,rst,matrix_A[11120],matrix_B[120],mul_res1[11120]);
multi_7x28 multi_7x28_mod_11121(clk,rst,matrix_A[11121],matrix_B[121],mul_res1[11121]);
multi_7x28 multi_7x28_mod_11122(clk,rst,matrix_A[11122],matrix_B[122],mul_res1[11122]);
multi_7x28 multi_7x28_mod_11123(clk,rst,matrix_A[11123],matrix_B[123],mul_res1[11123]);
multi_7x28 multi_7x28_mod_11124(clk,rst,matrix_A[11124],matrix_B[124],mul_res1[11124]);
multi_7x28 multi_7x28_mod_11125(clk,rst,matrix_A[11125],matrix_B[125],mul_res1[11125]);
multi_7x28 multi_7x28_mod_11126(clk,rst,matrix_A[11126],matrix_B[126],mul_res1[11126]);
multi_7x28 multi_7x28_mod_11127(clk,rst,matrix_A[11127],matrix_B[127],mul_res1[11127]);
multi_7x28 multi_7x28_mod_11128(clk,rst,matrix_A[11128],matrix_B[128],mul_res1[11128]);
multi_7x28 multi_7x28_mod_11129(clk,rst,matrix_A[11129],matrix_B[129],mul_res1[11129]);
multi_7x28 multi_7x28_mod_11130(clk,rst,matrix_A[11130],matrix_B[130],mul_res1[11130]);
multi_7x28 multi_7x28_mod_11131(clk,rst,matrix_A[11131],matrix_B[131],mul_res1[11131]);
multi_7x28 multi_7x28_mod_11132(clk,rst,matrix_A[11132],matrix_B[132],mul_res1[11132]);
multi_7x28 multi_7x28_mod_11133(clk,rst,matrix_A[11133],matrix_B[133],mul_res1[11133]);
multi_7x28 multi_7x28_mod_11134(clk,rst,matrix_A[11134],matrix_B[134],mul_res1[11134]);
multi_7x28 multi_7x28_mod_11135(clk,rst,matrix_A[11135],matrix_B[135],mul_res1[11135]);
multi_7x28 multi_7x28_mod_11136(clk,rst,matrix_A[11136],matrix_B[136],mul_res1[11136]);
multi_7x28 multi_7x28_mod_11137(clk,rst,matrix_A[11137],matrix_B[137],mul_res1[11137]);
multi_7x28 multi_7x28_mod_11138(clk,rst,matrix_A[11138],matrix_B[138],mul_res1[11138]);
multi_7x28 multi_7x28_mod_11139(clk,rst,matrix_A[11139],matrix_B[139],mul_res1[11139]);
multi_7x28 multi_7x28_mod_11140(clk,rst,matrix_A[11140],matrix_B[140],mul_res1[11140]);
multi_7x28 multi_7x28_mod_11141(clk,rst,matrix_A[11141],matrix_B[141],mul_res1[11141]);
multi_7x28 multi_7x28_mod_11142(clk,rst,matrix_A[11142],matrix_B[142],mul_res1[11142]);
multi_7x28 multi_7x28_mod_11143(clk,rst,matrix_A[11143],matrix_B[143],mul_res1[11143]);
multi_7x28 multi_7x28_mod_11144(clk,rst,matrix_A[11144],matrix_B[144],mul_res1[11144]);
multi_7x28 multi_7x28_mod_11145(clk,rst,matrix_A[11145],matrix_B[145],mul_res1[11145]);
multi_7x28 multi_7x28_mod_11146(clk,rst,matrix_A[11146],matrix_B[146],mul_res1[11146]);
multi_7x28 multi_7x28_mod_11147(clk,rst,matrix_A[11147],matrix_B[147],mul_res1[11147]);
multi_7x28 multi_7x28_mod_11148(clk,rst,matrix_A[11148],matrix_B[148],mul_res1[11148]);
multi_7x28 multi_7x28_mod_11149(clk,rst,matrix_A[11149],matrix_B[149],mul_res1[11149]);
multi_7x28 multi_7x28_mod_11150(clk,rst,matrix_A[11150],matrix_B[150],mul_res1[11150]);
multi_7x28 multi_7x28_mod_11151(clk,rst,matrix_A[11151],matrix_B[151],mul_res1[11151]);
multi_7x28 multi_7x28_mod_11152(clk,rst,matrix_A[11152],matrix_B[152],mul_res1[11152]);
multi_7x28 multi_7x28_mod_11153(clk,rst,matrix_A[11153],matrix_B[153],mul_res1[11153]);
multi_7x28 multi_7x28_mod_11154(clk,rst,matrix_A[11154],matrix_B[154],mul_res1[11154]);
multi_7x28 multi_7x28_mod_11155(clk,rst,matrix_A[11155],matrix_B[155],mul_res1[11155]);
multi_7x28 multi_7x28_mod_11156(clk,rst,matrix_A[11156],matrix_B[156],mul_res1[11156]);
multi_7x28 multi_7x28_mod_11157(clk,rst,matrix_A[11157],matrix_B[157],mul_res1[11157]);
multi_7x28 multi_7x28_mod_11158(clk,rst,matrix_A[11158],matrix_B[158],mul_res1[11158]);
multi_7x28 multi_7x28_mod_11159(clk,rst,matrix_A[11159],matrix_B[159],mul_res1[11159]);
multi_7x28 multi_7x28_mod_11160(clk,rst,matrix_A[11160],matrix_B[160],mul_res1[11160]);
multi_7x28 multi_7x28_mod_11161(clk,rst,matrix_A[11161],matrix_B[161],mul_res1[11161]);
multi_7x28 multi_7x28_mod_11162(clk,rst,matrix_A[11162],matrix_B[162],mul_res1[11162]);
multi_7x28 multi_7x28_mod_11163(clk,rst,matrix_A[11163],matrix_B[163],mul_res1[11163]);
multi_7x28 multi_7x28_mod_11164(clk,rst,matrix_A[11164],matrix_B[164],mul_res1[11164]);
multi_7x28 multi_7x28_mod_11165(clk,rst,matrix_A[11165],matrix_B[165],mul_res1[11165]);
multi_7x28 multi_7x28_mod_11166(clk,rst,matrix_A[11166],matrix_B[166],mul_res1[11166]);
multi_7x28 multi_7x28_mod_11167(clk,rst,matrix_A[11167],matrix_B[167],mul_res1[11167]);
multi_7x28 multi_7x28_mod_11168(clk,rst,matrix_A[11168],matrix_B[168],mul_res1[11168]);
multi_7x28 multi_7x28_mod_11169(clk,rst,matrix_A[11169],matrix_B[169],mul_res1[11169]);
multi_7x28 multi_7x28_mod_11170(clk,rst,matrix_A[11170],matrix_B[170],mul_res1[11170]);
multi_7x28 multi_7x28_mod_11171(clk,rst,matrix_A[11171],matrix_B[171],mul_res1[11171]);
multi_7x28 multi_7x28_mod_11172(clk,rst,matrix_A[11172],matrix_B[172],mul_res1[11172]);
multi_7x28 multi_7x28_mod_11173(clk,rst,matrix_A[11173],matrix_B[173],mul_res1[11173]);
multi_7x28 multi_7x28_mod_11174(clk,rst,matrix_A[11174],matrix_B[174],mul_res1[11174]);
multi_7x28 multi_7x28_mod_11175(clk,rst,matrix_A[11175],matrix_B[175],mul_res1[11175]);
multi_7x28 multi_7x28_mod_11176(clk,rst,matrix_A[11176],matrix_B[176],mul_res1[11176]);
multi_7x28 multi_7x28_mod_11177(clk,rst,matrix_A[11177],matrix_B[177],mul_res1[11177]);
multi_7x28 multi_7x28_mod_11178(clk,rst,matrix_A[11178],matrix_B[178],mul_res1[11178]);
multi_7x28 multi_7x28_mod_11179(clk,rst,matrix_A[11179],matrix_B[179],mul_res1[11179]);
multi_7x28 multi_7x28_mod_11180(clk,rst,matrix_A[11180],matrix_B[180],mul_res1[11180]);
multi_7x28 multi_7x28_mod_11181(clk,rst,matrix_A[11181],matrix_B[181],mul_res1[11181]);
multi_7x28 multi_7x28_mod_11182(clk,rst,matrix_A[11182],matrix_B[182],mul_res1[11182]);
multi_7x28 multi_7x28_mod_11183(clk,rst,matrix_A[11183],matrix_B[183],mul_res1[11183]);
multi_7x28 multi_7x28_mod_11184(clk,rst,matrix_A[11184],matrix_B[184],mul_res1[11184]);
multi_7x28 multi_7x28_mod_11185(clk,rst,matrix_A[11185],matrix_B[185],mul_res1[11185]);
multi_7x28 multi_7x28_mod_11186(clk,rst,matrix_A[11186],matrix_B[186],mul_res1[11186]);
multi_7x28 multi_7x28_mod_11187(clk,rst,matrix_A[11187],matrix_B[187],mul_res1[11187]);
multi_7x28 multi_7x28_mod_11188(clk,rst,matrix_A[11188],matrix_B[188],mul_res1[11188]);
multi_7x28 multi_7x28_mod_11189(clk,rst,matrix_A[11189],matrix_B[189],mul_res1[11189]);
multi_7x28 multi_7x28_mod_11190(clk,rst,matrix_A[11190],matrix_B[190],mul_res1[11190]);
multi_7x28 multi_7x28_mod_11191(clk,rst,matrix_A[11191],matrix_B[191],mul_res1[11191]);
multi_7x28 multi_7x28_mod_11192(clk,rst,matrix_A[11192],matrix_B[192],mul_res1[11192]);
multi_7x28 multi_7x28_mod_11193(clk,rst,matrix_A[11193],matrix_B[193],mul_res1[11193]);
multi_7x28 multi_7x28_mod_11194(clk,rst,matrix_A[11194],matrix_B[194],mul_res1[11194]);
multi_7x28 multi_7x28_mod_11195(clk,rst,matrix_A[11195],matrix_B[195],mul_res1[11195]);
multi_7x28 multi_7x28_mod_11196(clk,rst,matrix_A[11196],matrix_B[196],mul_res1[11196]);
multi_7x28 multi_7x28_mod_11197(clk,rst,matrix_A[11197],matrix_B[197],mul_res1[11197]);
multi_7x28 multi_7x28_mod_11198(clk,rst,matrix_A[11198],matrix_B[198],mul_res1[11198]);
multi_7x28 multi_7x28_mod_11199(clk,rst,matrix_A[11199],matrix_B[199],mul_res1[11199]);
multi_7x28 multi_7x28_mod_11200(clk,rst,matrix_A[11200],matrix_B[0],mul_res1[11200]);
multi_7x28 multi_7x28_mod_11201(clk,rst,matrix_A[11201],matrix_B[1],mul_res1[11201]);
multi_7x28 multi_7x28_mod_11202(clk,rst,matrix_A[11202],matrix_B[2],mul_res1[11202]);
multi_7x28 multi_7x28_mod_11203(clk,rst,matrix_A[11203],matrix_B[3],mul_res1[11203]);
multi_7x28 multi_7x28_mod_11204(clk,rst,matrix_A[11204],matrix_B[4],mul_res1[11204]);
multi_7x28 multi_7x28_mod_11205(clk,rst,matrix_A[11205],matrix_B[5],mul_res1[11205]);
multi_7x28 multi_7x28_mod_11206(clk,rst,matrix_A[11206],matrix_B[6],mul_res1[11206]);
multi_7x28 multi_7x28_mod_11207(clk,rst,matrix_A[11207],matrix_B[7],mul_res1[11207]);
multi_7x28 multi_7x28_mod_11208(clk,rst,matrix_A[11208],matrix_B[8],mul_res1[11208]);
multi_7x28 multi_7x28_mod_11209(clk,rst,matrix_A[11209],matrix_B[9],mul_res1[11209]);
multi_7x28 multi_7x28_mod_11210(clk,rst,matrix_A[11210],matrix_B[10],mul_res1[11210]);
multi_7x28 multi_7x28_mod_11211(clk,rst,matrix_A[11211],matrix_B[11],mul_res1[11211]);
multi_7x28 multi_7x28_mod_11212(clk,rst,matrix_A[11212],matrix_B[12],mul_res1[11212]);
multi_7x28 multi_7x28_mod_11213(clk,rst,matrix_A[11213],matrix_B[13],mul_res1[11213]);
multi_7x28 multi_7x28_mod_11214(clk,rst,matrix_A[11214],matrix_B[14],mul_res1[11214]);
multi_7x28 multi_7x28_mod_11215(clk,rst,matrix_A[11215],matrix_B[15],mul_res1[11215]);
multi_7x28 multi_7x28_mod_11216(clk,rst,matrix_A[11216],matrix_B[16],mul_res1[11216]);
multi_7x28 multi_7x28_mod_11217(clk,rst,matrix_A[11217],matrix_B[17],mul_res1[11217]);
multi_7x28 multi_7x28_mod_11218(clk,rst,matrix_A[11218],matrix_B[18],mul_res1[11218]);
multi_7x28 multi_7x28_mod_11219(clk,rst,matrix_A[11219],matrix_B[19],mul_res1[11219]);
multi_7x28 multi_7x28_mod_11220(clk,rst,matrix_A[11220],matrix_B[20],mul_res1[11220]);
multi_7x28 multi_7x28_mod_11221(clk,rst,matrix_A[11221],matrix_B[21],mul_res1[11221]);
multi_7x28 multi_7x28_mod_11222(clk,rst,matrix_A[11222],matrix_B[22],mul_res1[11222]);
multi_7x28 multi_7x28_mod_11223(clk,rst,matrix_A[11223],matrix_B[23],mul_res1[11223]);
multi_7x28 multi_7x28_mod_11224(clk,rst,matrix_A[11224],matrix_B[24],mul_res1[11224]);
multi_7x28 multi_7x28_mod_11225(clk,rst,matrix_A[11225],matrix_B[25],mul_res1[11225]);
multi_7x28 multi_7x28_mod_11226(clk,rst,matrix_A[11226],matrix_B[26],mul_res1[11226]);
multi_7x28 multi_7x28_mod_11227(clk,rst,matrix_A[11227],matrix_B[27],mul_res1[11227]);
multi_7x28 multi_7x28_mod_11228(clk,rst,matrix_A[11228],matrix_B[28],mul_res1[11228]);
multi_7x28 multi_7x28_mod_11229(clk,rst,matrix_A[11229],matrix_B[29],mul_res1[11229]);
multi_7x28 multi_7x28_mod_11230(clk,rst,matrix_A[11230],matrix_B[30],mul_res1[11230]);
multi_7x28 multi_7x28_mod_11231(clk,rst,matrix_A[11231],matrix_B[31],mul_res1[11231]);
multi_7x28 multi_7x28_mod_11232(clk,rst,matrix_A[11232],matrix_B[32],mul_res1[11232]);
multi_7x28 multi_7x28_mod_11233(clk,rst,matrix_A[11233],matrix_B[33],mul_res1[11233]);
multi_7x28 multi_7x28_mod_11234(clk,rst,matrix_A[11234],matrix_B[34],mul_res1[11234]);
multi_7x28 multi_7x28_mod_11235(clk,rst,matrix_A[11235],matrix_B[35],mul_res1[11235]);
multi_7x28 multi_7x28_mod_11236(clk,rst,matrix_A[11236],matrix_B[36],mul_res1[11236]);
multi_7x28 multi_7x28_mod_11237(clk,rst,matrix_A[11237],matrix_B[37],mul_res1[11237]);
multi_7x28 multi_7x28_mod_11238(clk,rst,matrix_A[11238],matrix_B[38],mul_res1[11238]);
multi_7x28 multi_7x28_mod_11239(clk,rst,matrix_A[11239],matrix_B[39],mul_res1[11239]);
multi_7x28 multi_7x28_mod_11240(clk,rst,matrix_A[11240],matrix_B[40],mul_res1[11240]);
multi_7x28 multi_7x28_mod_11241(clk,rst,matrix_A[11241],matrix_B[41],mul_res1[11241]);
multi_7x28 multi_7x28_mod_11242(clk,rst,matrix_A[11242],matrix_B[42],mul_res1[11242]);
multi_7x28 multi_7x28_mod_11243(clk,rst,matrix_A[11243],matrix_B[43],mul_res1[11243]);
multi_7x28 multi_7x28_mod_11244(clk,rst,matrix_A[11244],matrix_B[44],mul_res1[11244]);
multi_7x28 multi_7x28_mod_11245(clk,rst,matrix_A[11245],matrix_B[45],mul_res1[11245]);
multi_7x28 multi_7x28_mod_11246(clk,rst,matrix_A[11246],matrix_B[46],mul_res1[11246]);
multi_7x28 multi_7x28_mod_11247(clk,rst,matrix_A[11247],matrix_B[47],mul_res1[11247]);
multi_7x28 multi_7x28_mod_11248(clk,rst,matrix_A[11248],matrix_B[48],mul_res1[11248]);
multi_7x28 multi_7x28_mod_11249(clk,rst,matrix_A[11249],matrix_B[49],mul_res1[11249]);
multi_7x28 multi_7x28_mod_11250(clk,rst,matrix_A[11250],matrix_B[50],mul_res1[11250]);
multi_7x28 multi_7x28_mod_11251(clk,rst,matrix_A[11251],matrix_B[51],mul_res1[11251]);
multi_7x28 multi_7x28_mod_11252(clk,rst,matrix_A[11252],matrix_B[52],mul_res1[11252]);
multi_7x28 multi_7x28_mod_11253(clk,rst,matrix_A[11253],matrix_B[53],mul_res1[11253]);
multi_7x28 multi_7x28_mod_11254(clk,rst,matrix_A[11254],matrix_B[54],mul_res1[11254]);
multi_7x28 multi_7x28_mod_11255(clk,rst,matrix_A[11255],matrix_B[55],mul_res1[11255]);
multi_7x28 multi_7x28_mod_11256(clk,rst,matrix_A[11256],matrix_B[56],mul_res1[11256]);
multi_7x28 multi_7x28_mod_11257(clk,rst,matrix_A[11257],matrix_B[57],mul_res1[11257]);
multi_7x28 multi_7x28_mod_11258(clk,rst,matrix_A[11258],matrix_B[58],mul_res1[11258]);
multi_7x28 multi_7x28_mod_11259(clk,rst,matrix_A[11259],matrix_B[59],mul_res1[11259]);
multi_7x28 multi_7x28_mod_11260(clk,rst,matrix_A[11260],matrix_B[60],mul_res1[11260]);
multi_7x28 multi_7x28_mod_11261(clk,rst,matrix_A[11261],matrix_B[61],mul_res1[11261]);
multi_7x28 multi_7x28_mod_11262(clk,rst,matrix_A[11262],matrix_B[62],mul_res1[11262]);
multi_7x28 multi_7x28_mod_11263(clk,rst,matrix_A[11263],matrix_B[63],mul_res1[11263]);
multi_7x28 multi_7x28_mod_11264(clk,rst,matrix_A[11264],matrix_B[64],mul_res1[11264]);
multi_7x28 multi_7x28_mod_11265(clk,rst,matrix_A[11265],matrix_B[65],mul_res1[11265]);
multi_7x28 multi_7x28_mod_11266(clk,rst,matrix_A[11266],matrix_B[66],mul_res1[11266]);
multi_7x28 multi_7x28_mod_11267(clk,rst,matrix_A[11267],matrix_B[67],mul_res1[11267]);
multi_7x28 multi_7x28_mod_11268(clk,rst,matrix_A[11268],matrix_B[68],mul_res1[11268]);
multi_7x28 multi_7x28_mod_11269(clk,rst,matrix_A[11269],matrix_B[69],mul_res1[11269]);
multi_7x28 multi_7x28_mod_11270(clk,rst,matrix_A[11270],matrix_B[70],mul_res1[11270]);
multi_7x28 multi_7x28_mod_11271(clk,rst,matrix_A[11271],matrix_B[71],mul_res1[11271]);
multi_7x28 multi_7x28_mod_11272(clk,rst,matrix_A[11272],matrix_B[72],mul_res1[11272]);
multi_7x28 multi_7x28_mod_11273(clk,rst,matrix_A[11273],matrix_B[73],mul_res1[11273]);
multi_7x28 multi_7x28_mod_11274(clk,rst,matrix_A[11274],matrix_B[74],mul_res1[11274]);
multi_7x28 multi_7x28_mod_11275(clk,rst,matrix_A[11275],matrix_B[75],mul_res1[11275]);
multi_7x28 multi_7x28_mod_11276(clk,rst,matrix_A[11276],matrix_B[76],mul_res1[11276]);
multi_7x28 multi_7x28_mod_11277(clk,rst,matrix_A[11277],matrix_B[77],mul_res1[11277]);
multi_7x28 multi_7x28_mod_11278(clk,rst,matrix_A[11278],matrix_B[78],mul_res1[11278]);
multi_7x28 multi_7x28_mod_11279(clk,rst,matrix_A[11279],matrix_B[79],mul_res1[11279]);
multi_7x28 multi_7x28_mod_11280(clk,rst,matrix_A[11280],matrix_B[80],mul_res1[11280]);
multi_7x28 multi_7x28_mod_11281(clk,rst,matrix_A[11281],matrix_B[81],mul_res1[11281]);
multi_7x28 multi_7x28_mod_11282(clk,rst,matrix_A[11282],matrix_B[82],mul_res1[11282]);
multi_7x28 multi_7x28_mod_11283(clk,rst,matrix_A[11283],matrix_B[83],mul_res1[11283]);
multi_7x28 multi_7x28_mod_11284(clk,rst,matrix_A[11284],matrix_B[84],mul_res1[11284]);
multi_7x28 multi_7x28_mod_11285(clk,rst,matrix_A[11285],matrix_B[85],mul_res1[11285]);
multi_7x28 multi_7x28_mod_11286(clk,rst,matrix_A[11286],matrix_B[86],mul_res1[11286]);
multi_7x28 multi_7x28_mod_11287(clk,rst,matrix_A[11287],matrix_B[87],mul_res1[11287]);
multi_7x28 multi_7x28_mod_11288(clk,rst,matrix_A[11288],matrix_B[88],mul_res1[11288]);
multi_7x28 multi_7x28_mod_11289(clk,rst,matrix_A[11289],matrix_B[89],mul_res1[11289]);
multi_7x28 multi_7x28_mod_11290(clk,rst,matrix_A[11290],matrix_B[90],mul_res1[11290]);
multi_7x28 multi_7x28_mod_11291(clk,rst,matrix_A[11291],matrix_B[91],mul_res1[11291]);
multi_7x28 multi_7x28_mod_11292(clk,rst,matrix_A[11292],matrix_B[92],mul_res1[11292]);
multi_7x28 multi_7x28_mod_11293(clk,rst,matrix_A[11293],matrix_B[93],mul_res1[11293]);
multi_7x28 multi_7x28_mod_11294(clk,rst,matrix_A[11294],matrix_B[94],mul_res1[11294]);
multi_7x28 multi_7x28_mod_11295(clk,rst,matrix_A[11295],matrix_B[95],mul_res1[11295]);
multi_7x28 multi_7x28_mod_11296(clk,rst,matrix_A[11296],matrix_B[96],mul_res1[11296]);
multi_7x28 multi_7x28_mod_11297(clk,rst,matrix_A[11297],matrix_B[97],mul_res1[11297]);
multi_7x28 multi_7x28_mod_11298(clk,rst,matrix_A[11298],matrix_B[98],mul_res1[11298]);
multi_7x28 multi_7x28_mod_11299(clk,rst,matrix_A[11299],matrix_B[99],mul_res1[11299]);
multi_7x28 multi_7x28_mod_11300(clk,rst,matrix_A[11300],matrix_B[100],mul_res1[11300]);
multi_7x28 multi_7x28_mod_11301(clk,rst,matrix_A[11301],matrix_B[101],mul_res1[11301]);
multi_7x28 multi_7x28_mod_11302(clk,rst,matrix_A[11302],matrix_B[102],mul_res1[11302]);
multi_7x28 multi_7x28_mod_11303(clk,rst,matrix_A[11303],matrix_B[103],mul_res1[11303]);
multi_7x28 multi_7x28_mod_11304(clk,rst,matrix_A[11304],matrix_B[104],mul_res1[11304]);
multi_7x28 multi_7x28_mod_11305(clk,rst,matrix_A[11305],matrix_B[105],mul_res1[11305]);
multi_7x28 multi_7x28_mod_11306(clk,rst,matrix_A[11306],matrix_B[106],mul_res1[11306]);
multi_7x28 multi_7x28_mod_11307(clk,rst,matrix_A[11307],matrix_B[107],mul_res1[11307]);
multi_7x28 multi_7x28_mod_11308(clk,rst,matrix_A[11308],matrix_B[108],mul_res1[11308]);
multi_7x28 multi_7x28_mod_11309(clk,rst,matrix_A[11309],matrix_B[109],mul_res1[11309]);
multi_7x28 multi_7x28_mod_11310(clk,rst,matrix_A[11310],matrix_B[110],mul_res1[11310]);
multi_7x28 multi_7x28_mod_11311(clk,rst,matrix_A[11311],matrix_B[111],mul_res1[11311]);
multi_7x28 multi_7x28_mod_11312(clk,rst,matrix_A[11312],matrix_B[112],mul_res1[11312]);
multi_7x28 multi_7x28_mod_11313(clk,rst,matrix_A[11313],matrix_B[113],mul_res1[11313]);
multi_7x28 multi_7x28_mod_11314(clk,rst,matrix_A[11314],matrix_B[114],mul_res1[11314]);
multi_7x28 multi_7x28_mod_11315(clk,rst,matrix_A[11315],matrix_B[115],mul_res1[11315]);
multi_7x28 multi_7x28_mod_11316(clk,rst,matrix_A[11316],matrix_B[116],mul_res1[11316]);
multi_7x28 multi_7x28_mod_11317(clk,rst,matrix_A[11317],matrix_B[117],mul_res1[11317]);
multi_7x28 multi_7x28_mod_11318(clk,rst,matrix_A[11318],matrix_B[118],mul_res1[11318]);
multi_7x28 multi_7x28_mod_11319(clk,rst,matrix_A[11319],matrix_B[119],mul_res1[11319]);
multi_7x28 multi_7x28_mod_11320(clk,rst,matrix_A[11320],matrix_B[120],mul_res1[11320]);
multi_7x28 multi_7x28_mod_11321(clk,rst,matrix_A[11321],matrix_B[121],mul_res1[11321]);
multi_7x28 multi_7x28_mod_11322(clk,rst,matrix_A[11322],matrix_B[122],mul_res1[11322]);
multi_7x28 multi_7x28_mod_11323(clk,rst,matrix_A[11323],matrix_B[123],mul_res1[11323]);
multi_7x28 multi_7x28_mod_11324(clk,rst,matrix_A[11324],matrix_B[124],mul_res1[11324]);
multi_7x28 multi_7x28_mod_11325(clk,rst,matrix_A[11325],matrix_B[125],mul_res1[11325]);
multi_7x28 multi_7x28_mod_11326(clk,rst,matrix_A[11326],matrix_B[126],mul_res1[11326]);
multi_7x28 multi_7x28_mod_11327(clk,rst,matrix_A[11327],matrix_B[127],mul_res1[11327]);
multi_7x28 multi_7x28_mod_11328(clk,rst,matrix_A[11328],matrix_B[128],mul_res1[11328]);
multi_7x28 multi_7x28_mod_11329(clk,rst,matrix_A[11329],matrix_B[129],mul_res1[11329]);
multi_7x28 multi_7x28_mod_11330(clk,rst,matrix_A[11330],matrix_B[130],mul_res1[11330]);
multi_7x28 multi_7x28_mod_11331(clk,rst,matrix_A[11331],matrix_B[131],mul_res1[11331]);
multi_7x28 multi_7x28_mod_11332(clk,rst,matrix_A[11332],matrix_B[132],mul_res1[11332]);
multi_7x28 multi_7x28_mod_11333(clk,rst,matrix_A[11333],matrix_B[133],mul_res1[11333]);
multi_7x28 multi_7x28_mod_11334(clk,rst,matrix_A[11334],matrix_B[134],mul_res1[11334]);
multi_7x28 multi_7x28_mod_11335(clk,rst,matrix_A[11335],matrix_B[135],mul_res1[11335]);
multi_7x28 multi_7x28_mod_11336(clk,rst,matrix_A[11336],matrix_B[136],mul_res1[11336]);
multi_7x28 multi_7x28_mod_11337(clk,rst,matrix_A[11337],matrix_B[137],mul_res1[11337]);
multi_7x28 multi_7x28_mod_11338(clk,rst,matrix_A[11338],matrix_B[138],mul_res1[11338]);
multi_7x28 multi_7x28_mod_11339(clk,rst,matrix_A[11339],matrix_B[139],mul_res1[11339]);
multi_7x28 multi_7x28_mod_11340(clk,rst,matrix_A[11340],matrix_B[140],mul_res1[11340]);
multi_7x28 multi_7x28_mod_11341(clk,rst,matrix_A[11341],matrix_B[141],mul_res1[11341]);
multi_7x28 multi_7x28_mod_11342(clk,rst,matrix_A[11342],matrix_B[142],mul_res1[11342]);
multi_7x28 multi_7x28_mod_11343(clk,rst,matrix_A[11343],matrix_B[143],mul_res1[11343]);
multi_7x28 multi_7x28_mod_11344(clk,rst,matrix_A[11344],matrix_B[144],mul_res1[11344]);
multi_7x28 multi_7x28_mod_11345(clk,rst,matrix_A[11345],matrix_B[145],mul_res1[11345]);
multi_7x28 multi_7x28_mod_11346(clk,rst,matrix_A[11346],matrix_B[146],mul_res1[11346]);
multi_7x28 multi_7x28_mod_11347(clk,rst,matrix_A[11347],matrix_B[147],mul_res1[11347]);
multi_7x28 multi_7x28_mod_11348(clk,rst,matrix_A[11348],matrix_B[148],mul_res1[11348]);
multi_7x28 multi_7x28_mod_11349(clk,rst,matrix_A[11349],matrix_B[149],mul_res1[11349]);
multi_7x28 multi_7x28_mod_11350(clk,rst,matrix_A[11350],matrix_B[150],mul_res1[11350]);
multi_7x28 multi_7x28_mod_11351(clk,rst,matrix_A[11351],matrix_B[151],mul_res1[11351]);
multi_7x28 multi_7x28_mod_11352(clk,rst,matrix_A[11352],matrix_B[152],mul_res1[11352]);
multi_7x28 multi_7x28_mod_11353(clk,rst,matrix_A[11353],matrix_B[153],mul_res1[11353]);
multi_7x28 multi_7x28_mod_11354(clk,rst,matrix_A[11354],matrix_B[154],mul_res1[11354]);
multi_7x28 multi_7x28_mod_11355(clk,rst,matrix_A[11355],matrix_B[155],mul_res1[11355]);
multi_7x28 multi_7x28_mod_11356(clk,rst,matrix_A[11356],matrix_B[156],mul_res1[11356]);
multi_7x28 multi_7x28_mod_11357(clk,rst,matrix_A[11357],matrix_B[157],mul_res1[11357]);
multi_7x28 multi_7x28_mod_11358(clk,rst,matrix_A[11358],matrix_B[158],mul_res1[11358]);
multi_7x28 multi_7x28_mod_11359(clk,rst,matrix_A[11359],matrix_B[159],mul_res1[11359]);
multi_7x28 multi_7x28_mod_11360(clk,rst,matrix_A[11360],matrix_B[160],mul_res1[11360]);
multi_7x28 multi_7x28_mod_11361(clk,rst,matrix_A[11361],matrix_B[161],mul_res1[11361]);
multi_7x28 multi_7x28_mod_11362(clk,rst,matrix_A[11362],matrix_B[162],mul_res1[11362]);
multi_7x28 multi_7x28_mod_11363(clk,rst,matrix_A[11363],matrix_B[163],mul_res1[11363]);
multi_7x28 multi_7x28_mod_11364(clk,rst,matrix_A[11364],matrix_B[164],mul_res1[11364]);
multi_7x28 multi_7x28_mod_11365(clk,rst,matrix_A[11365],matrix_B[165],mul_res1[11365]);
multi_7x28 multi_7x28_mod_11366(clk,rst,matrix_A[11366],matrix_B[166],mul_res1[11366]);
multi_7x28 multi_7x28_mod_11367(clk,rst,matrix_A[11367],matrix_B[167],mul_res1[11367]);
multi_7x28 multi_7x28_mod_11368(clk,rst,matrix_A[11368],matrix_B[168],mul_res1[11368]);
multi_7x28 multi_7x28_mod_11369(clk,rst,matrix_A[11369],matrix_B[169],mul_res1[11369]);
multi_7x28 multi_7x28_mod_11370(clk,rst,matrix_A[11370],matrix_B[170],mul_res1[11370]);
multi_7x28 multi_7x28_mod_11371(clk,rst,matrix_A[11371],matrix_B[171],mul_res1[11371]);
multi_7x28 multi_7x28_mod_11372(clk,rst,matrix_A[11372],matrix_B[172],mul_res1[11372]);
multi_7x28 multi_7x28_mod_11373(clk,rst,matrix_A[11373],matrix_B[173],mul_res1[11373]);
multi_7x28 multi_7x28_mod_11374(clk,rst,matrix_A[11374],matrix_B[174],mul_res1[11374]);
multi_7x28 multi_7x28_mod_11375(clk,rst,matrix_A[11375],matrix_B[175],mul_res1[11375]);
multi_7x28 multi_7x28_mod_11376(clk,rst,matrix_A[11376],matrix_B[176],mul_res1[11376]);
multi_7x28 multi_7x28_mod_11377(clk,rst,matrix_A[11377],matrix_B[177],mul_res1[11377]);
multi_7x28 multi_7x28_mod_11378(clk,rst,matrix_A[11378],matrix_B[178],mul_res1[11378]);
multi_7x28 multi_7x28_mod_11379(clk,rst,matrix_A[11379],matrix_B[179],mul_res1[11379]);
multi_7x28 multi_7x28_mod_11380(clk,rst,matrix_A[11380],matrix_B[180],mul_res1[11380]);
multi_7x28 multi_7x28_mod_11381(clk,rst,matrix_A[11381],matrix_B[181],mul_res1[11381]);
multi_7x28 multi_7x28_mod_11382(clk,rst,matrix_A[11382],matrix_B[182],mul_res1[11382]);
multi_7x28 multi_7x28_mod_11383(clk,rst,matrix_A[11383],matrix_B[183],mul_res1[11383]);
multi_7x28 multi_7x28_mod_11384(clk,rst,matrix_A[11384],matrix_B[184],mul_res1[11384]);
multi_7x28 multi_7x28_mod_11385(clk,rst,matrix_A[11385],matrix_B[185],mul_res1[11385]);
multi_7x28 multi_7x28_mod_11386(clk,rst,matrix_A[11386],matrix_B[186],mul_res1[11386]);
multi_7x28 multi_7x28_mod_11387(clk,rst,matrix_A[11387],matrix_B[187],mul_res1[11387]);
multi_7x28 multi_7x28_mod_11388(clk,rst,matrix_A[11388],matrix_B[188],mul_res1[11388]);
multi_7x28 multi_7x28_mod_11389(clk,rst,matrix_A[11389],matrix_B[189],mul_res1[11389]);
multi_7x28 multi_7x28_mod_11390(clk,rst,matrix_A[11390],matrix_B[190],mul_res1[11390]);
multi_7x28 multi_7x28_mod_11391(clk,rst,matrix_A[11391],matrix_B[191],mul_res1[11391]);
multi_7x28 multi_7x28_mod_11392(clk,rst,matrix_A[11392],matrix_B[192],mul_res1[11392]);
multi_7x28 multi_7x28_mod_11393(clk,rst,matrix_A[11393],matrix_B[193],mul_res1[11393]);
multi_7x28 multi_7x28_mod_11394(clk,rst,matrix_A[11394],matrix_B[194],mul_res1[11394]);
multi_7x28 multi_7x28_mod_11395(clk,rst,matrix_A[11395],matrix_B[195],mul_res1[11395]);
multi_7x28 multi_7x28_mod_11396(clk,rst,matrix_A[11396],matrix_B[196],mul_res1[11396]);
multi_7x28 multi_7x28_mod_11397(clk,rst,matrix_A[11397],matrix_B[197],mul_res1[11397]);
multi_7x28 multi_7x28_mod_11398(clk,rst,matrix_A[11398],matrix_B[198],mul_res1[11398]);
multi_7x28 multi_7x28_mod_11399(clk,rst,matrix_A[11399],matrix_B[199],mul_res1[11399]);
multi_7x28 multi_7x28_mod_11400(clk,rst,matrix_A[11400],matrix_B[0],mul_res1[11400]);
multi_7x28 multi_7x28_mod_11401(clk,rst,matrix_A[11401],matrix_B[1],mul_res1[11401]);
multi_7x28 multi_7x28_mod_11402(clk,rst,matrix_A[11402],matrix_B[2],mul_res1[11402]);
multi_7x28 multi_7x28_mod_11403(clk,rst,matrix_A[11403],matrix_B[3],mul_res1[11403]);
multi_7x28 multi_7x28_mod_11404(clk,rst,matrix_A[11404],matrix_B[4],mul_res1[11404]);
multi_7x28 multi_7x28_mod_11405(clk,rst,matrix_A[11405],matrix_B[5],mul_res1[11405]);
multi_7x28 multi_7x28_mod_11406(clk,rst,matrix_A[11406],matrix_B[6],mul_res1[11406]);
multi_7x28 multi_7x28_mod_11407(clk,rst,matrix_A[11407],matrix_B[7],mul_res1[11407]);
multi_7x28 multi_7x28_mod_11408(clk,rst,matrix_A[11408],matrix_B[8],mul_res1[11408]);
multi_7x28 multi_7x28_mod_11409(clk,rst,matrix_A[11409],matrix_B[9],mul_res1[11409]);
multi_7x28 multi_7x28_mod_11410(clk,rst,matrix_A[11410],matrix_B[10],mul_res1[11410]);
multi_7x28 multi_7x28_mod_11411(clk,rst,matrix_A[11411],matrix_B[11],mul_res1[11411]);
multi_7x28 multi_7x28_mod_11412(clk,rst,matrix_A[11412],matrix_B[12],mul_res1[11412]);
multi_7x28 multi_7x28_mod_11413(clk,rst,matrix_A[11413],matrix_B[13],mul_res1[11413]);
multi_7x28 multi_7x28_mod_11414(clk,rst,matrix_A[11414],matrix_B[14],mul_res1[11414]);
multi_7x28 multi_7x28_mod_11415(clk,rst,matrix_A[11415],matrix_B[15],mul_res1[11415]);
multi_7x28 multi_7x28_mod_11416(clk,rst,matrix_A[11416],matrix_B[16],mul_res1[11416]);
multi_7x28 multi_7x28_mod_11417(clk,rst,matrix_A[11417],matrix_B[17],mul_res1[11417]);
multi_7x28 multi_7x28_mod_11418(clk,rst,matrix_A[11418],matrix_B[18],mul_res1[11418]);
multi_7x28 multi_7x28_mod_11419(clk,rst,matrix_A[11419],matrix_B[19],mul_res1[11419]);
multi_7x28 multi_7x28_mod_11420(clk,rst,matrix_A[11420],matrix_B[20],mul_res1[11420]);
multi_7x28 multi_7x28_mod_11421(clk,rst,matrix_A[11421],matrix_B[21],mul_res1[11421]);
multi_7x28 multi_7x28_mod_11422(clk,rst,matrix_A[11422],matrix_B[22],mul_res1[11422]);
multi_7x28 multi_7x28_mod_11423(clk,rst,matrix_A[11423],matrix_B[23],mul_res1[11423]);
multi_7x28 multi_7x28_mod_11424(clk,rst,matrix_A[11424],matrix_B[24],mul_res1[11424]);
multi_7x28 multi_7x28_mod_11425(clk,rst,matrix_A[11425],matrix_B[25],mul_res1[11425]);
multi_7x28 multi_7x28_mod_11426(clk,rst,matrix_A[11426],matrix_B[26],mul_res1[11426]);
multi_7x28 multi_7x28_mod_11427(clk,rst,matrix_A[11427],matrix_B[27],mul_res1[11427]);
multi_7x28 multi_7x28_mod_11428(clk,rst,matrix_A[11428],matrix_B[28],mul_res1[11428]);
multi_7x28 multi_7x28_mod_11429(clk,rst,matrix_A[11429],matrix_B[29],mul_res1[11429]);
multi_7x28 multi_7x28_mod_11430(clk,rst,matrix_A[11430],matrix_B[30],mul_res1[11430]);
multi_7x28 multi_7x28_mod_11431(clk,rst,matrix_A[11431],matrix_B[31],mul_res1[11431]);
multi_7x28 multi_7x28_mod_11432(clk,rst,matrix_A[11432],matrix_B[32],mul_res1[11432]);
multi_7x28 multi_7x28_mod_11433(clk,rst,matrix_A[11433],matrix_B[33],mul_res1[11433]);
multi_7x28 multi_7x28_mod_11434(clk,rst,matrix_A[11434],matrix_B[34],mul_res1[11434]);
multi_7x28 multi_7x28_mod_11435(clk,rst,matrix_A[11435],matrix_B[35],mul_res1[11435]);
multi_7x28 multi_7x28_mod_11436(clk,rst,matrix_A[11436],matrix_B[36],mul_res1[11436]);
multi_7x28 multi_7x28_mod_11437(clk,rst,matrix_A[11437],matrix_B[37],mul_res1[11437]);
multi_7x28 multi_7x28_mod_11438(clk,rst,matrix_A[11438],matrix_B[38],mul_res1[11438]);
multi_7x28 multi_7x28_mod_11439(clk,rst,matrix_A[11439],matrix_B[39],mul_res1[11439]);
multi_7x28 multi_7x28_mod_11440(clk,rst,matrix_A[11440],matrix_B[40],mul_res1[11440]);
multi_7x28 multi_7x28_mod_11441(clk,rst,matrix_A[11441],matrix_B[41],mul_res1[11441]);
multi_7x28 multi_7x28_mod_11442(clk,rst,matrix_A[11442],matrix_B[42],mul_res1[11442]);
multi_7x28 multi_7x28_mod_11443(clk,rst,matrix_A[11443],matrix_B[43],mul_res1[11443]);
multi_7x28 multi_7x28_mod_11444(clk,rst,matrix_A[11444],matrix_B[44],mul_res1[11444]);
multi_7x28 multi_7x28_mod_11445(clk,rst,matrix_A[11445],matrix_B[45],mul_res1[11445]);
multi_7x28 multi_7x28_mod_11446(clk,rst,matrix_A[11446],matrix_B[46],mul_res1[11446]);
multi_7x28 multi_7x28_mod_11447(clk,rst,matrix_A[11447],matrix_B[47],mul_res1[11447]);
multi_7x28 multi_7x28_mod_11448(clk,rst,matrix_A[11448],matrix_B[48],mul_res1[11448]);
multi_7x28 multi_7x28_mod_11449(clk,rst,matrix_A[11449],matrix_B[49],mul_res1[11449]);
multi_7x28 multi_7x28_mod_11450(clk,rst,matrix_A[11450],matrix_B[50],mul_res1[11450]);
multi_7x28 multi_7x28_mod_11451(clk,rst,matrix_A[11451],matrix_B[51],mul_res1[11451]);
multi_7x28 multi_7x28_mod_11452(clk,rst,matrix_A[11452],matrix_B[52],mul_res1[11452]);
multi_7x28 multi_7x28_mod_11453(clk,rst,matrix_A[11453],matrix_B[53],mul_res1[11453]);
multi_7x28 multi_7x28_mod_11454(clk,rst,matrix_A[11454],matrix_B[54],mul_res1[11454]);
multi_7x28 multi_7x28_mod_11455(clk,rst,matrix_A[11455],matrix_B[55],mul_res1[11455]);
multi_7x28 multi_7x28_mod_11456(clk,rst,matrix_A[11456],matrix_B[56],mul_res1[11456]);
multi_7x28 multi_7x28_mod_11457(clk,rst,matrix_A[11457],matrix_B[57],mul_res1[11457]);
multi_7x28 multi_7x28_mod_11458(clk,rst,matrix_A[11458],matrix_B[58],mul_res1[11458]);
multi_7x28 multi_7x28_mod_11459(clk,rst,matrix_A[11459],matrix_B[59],mul_res1[11459]);
multi_7x28 multi_7x28_mod_11460(clk,rst,matrix_A[11460],matrix_B[60],mul_res1[11460]);
multi_7x28 multi_7x28_mod_11461(clk,rst,matrix_A[11461],matrix_B[61],mul_res1[11461]);
multi_7x28 multi_7x28_mod_11462(clk,rst,matrix_A[11462],matrix_B[62],mul_res1[11462]);
multi_7x28 multi_7x28_mod_11463(clk,rst,matrix_A[11463],matrix_B[63],mul_res1[11463]);
multi_7x28 multi_7x28_mod_11464(clk,rst,matrix_A[11464],matrix_B[64],mul_res1[11464]);
multi_7x28 multi_7x28_mod_11465(clk,rst,matrix_A[11465],matrix_B[65],mul_res1[11465]);
multi_7x28 multi_7x28_mod_11466(clk,rst,matrix_A[11466],matrix_B[66],mul_res1[11466]);
multi_7x28 multi_7x28_mod_11467(clk,rst,matrix_A[11467],matrix_B[67],mul_res1[11467]);
multi_7x28 multi_7x28_mod_11468(clk,rst,matrix_A[11468],matrix_B[68],mul_res1[11468]);
multi_7x28 multi_7x28_mod_11469(clk,rst,matrix_A[11469],matrix_B[69],mul_res1[11469]);
multi_7x28 multi_7x28_mod_11470(clk,rst,matrix_A[11470],matrix_B[70],mul_res1[11470]);
multi_7x28 multi_7x28_mod_11471(clk,rst,matrix_A[11471],matrix_B[71],mul_res1[11471]);
multi_7x28 multi_7x28_mod_11472(clk,rst,matrix_A[11472],matrix_B[72],mul_res1[11472]);
multi_7x28 multi_7x28_mod_11473(clk,rst,matrix_A[11473],matrix_B[73],mul_res1[11473]);
multi_7x28 multi_7x28_mod_11474(clk,rst,matrix_A[11474],matrix_B[74],mul_res1[11474]);
multi_7x28 multi_7x28_mod_11475(clk,rst,matrix_A[11475],matrix_B[75],mul_res1[11475]);
multi_7x28 multi_7x28_mod_11476(clk,rst,matrix_A[11476],matrix_B[76],mul_res1[11476]);
multi_7x28 multi_7x28_mod_11477(clk,rst,matrix_A[11477],matrix_B[77],mul_res1[11477]);
multi_7x28 multi_7x28_mod_11478(clk,rst,matrix_A[11478],matrix_B[78],mul_res1[11478]);
multi_7x28 multi_7x28_mod_11479(clk,rst,matrix_A[11479],matrix_B[79],mul_res1[11479]);
multi_7x28 multi_7x28_mod_11480(clk,rst,matrix_A[11480],matrix_B[80],mul_res1[11480]);
multi_7x28 multi_7x28_mod_11481(clk,rst,matrix_A[11481],matrix_B[81],mul_res1[11481]);
multi_7x28 multi_7x28_mod_11482(clk,rst,matrix_A[11482],matrix_B[82],mul_res1[11482]);
multi_7x28 multi_7x28_mod_11483(clk,rst,matrix_A[11483],matrix_B[83],mul_res1[11483]);
multi_7x28 multi_7x28_mod_11484(clk,rst,matrix_A[11484],matrix_B[84],mul_res1[11484]);
multi_7x28 multi_7x28_mod_11485(clk,rst,matrix_A[11485],matrix_B[85],mul_res1[11485]);
multi_7x28 multi_7x28_mod_11486(clk,rst,matrix_A[11486],matrix_B[86],mul_res1[11486]);
multi_7x28 multi_7x28_mod_11487(clk,rst,matrix_A[11487],matrix_B[87],mul_res1[11487]);
multi_7x28 multi_7x28_mod_11488(clk,rst,matrix_A[11488],matrix_B[88],mul_res1[11488]);
multi_7x28 multi_7x28_mod_11489(clk,rst,matrix_A[11489],matrix_B[89],mul_res1[11489]);
multi_7x28 multi_7x28_mod_11490(clk,rst,matrix_A[11490],matrix_B[90],mul_res1[11490]);
multi_7x28 multi_7x28_mod_11491(clk,rst,matrix_A[11491],matrix_B[91],mul_res1[11491]);
multi_7x28 multi_7x28_mod_11492(clk,rst,matrix_A[11492],matrix_B[92],mul_res1[11492]);
multi_7x28 multi_7x28_mod_11493(clk,rst,matrix_A[11493],matrix_B[93],mul_res1[11493]);
multi_7x28 multi_7x28_mod_11494(clk,rst,matrix_A[11494],matrix_B[94],mul_res1[11494]);
multi_7x28 multi_7x28_mod_11495(clk,rst,matrix_A[11495],matrix_B[95],mul_res1[11495]);
multi_7x28 multi_7x28_mod_11496(clk,rst,matrix_A[11496],matrix_B[96],mul_res1[11496]);
multi_7x28 multi_7x28_mod_11497(clk,rst,matrix_A[11497],matrix_B[97],mul_res1[11497]);
multi_7x28 multi_7x28_mod_11498(clk,rst,matrix_A[11498],matrix_B[98],mul_res1[11498]);
multi_7x28 multi_7x28_mod_11499(clk,rst,matrix_A[11499],matrix_B[99],mul_res1[11499]);
multi_7x28 multi_7x28_mod_11500(clk,rst,matrix_A[11500],matrix_B[100],mul_res1[11500]);
multi_7x28 multi_7x28_mod_11501(clk,rst,matrix_A[11501],matrix_B[101],mul_res1[11501]);
multi_7x28 multi_7x28_mod_11502(clk,rst,matrix_A[11502],matrix_B[102],mul_res1[11502]);
multi_7x28 multi_7x28_mod_11503(clk,rst,matrix_A[11503],matrix_B[103],mul_res1[11503]);
multi_7x28 multi_7x28_mod_11504(clk,rst,matrix_A[11504],matrix_B[104],mul_res1[11504]);
multi_7x28 multi_7x28_mod_11505(clk,rst,matrix_A[11505],matrix_B[105],mul_res1[11505]);
multi_7x28 multi_7x28_mod_11506(clk,rst,matrix_A[11506],matrix_B[106],mul_res1[11506]);
multi_7x28 multi_7x28_mod_11507(clk,rst,matrix_A[11507],matrix_B[107],mul_res1[11507]);
multi_7x28 multi_7x28_mod_11508(clk,rst,matrix_A[11508],matrix_B[108],mul_res1[11508]);
multi_7x28 multi_7x28_mod_11509(clk,rst,matrix_A[11509],matrix_B[109],mul_res1[11509]);
multi_7x28 multi_7x28_mod_11510(clk,rst,matrix_A[11510],matrix_B[110],mul_res1[11510]);
multi_7x28 multi_7x28_mod_11511(clk,rst,matrix_A[11511],matrix_B[111],mul_res1[11511]);
multi_7x28 multi_7x28_mod_11512(clk,rst,matrix_A[11512],matrix_B[112],mul_res1[11512]);
multi_7x28 multi_7x28_mod_11513(clk,rst,matrix_A[11513],matrix_B[113],mul_res1[11513]);
multi_7x28 multi_7x28_mod_11514(clk,rst,matrix_A[11514],matrix_B[114],mul_res1[11514]);
multi_7x28 multi_7x28_mod_11515(clk,rst,matrix_A[11515],matrix_B[115],mul_res1[11515]);
multi_7x28 multi_7x28_mod_11516(clk,rst,matrix_A[11516],matrix_B[116],mul_res1[11516]);
multi_7x28 multi_7x28_mod_11517(clk,rst,matrix_A[11517],matrix_B[117],mul_res1[11517]);
multi_7x28 multi_7x28_mod_11518(clk,rst,matrix_A[11518],matrix_B[118],mul_res1[11518]);
multi_7x28 multi_7x28_mod_11519(clk,rst,matrix_A[11519],matrix_B[119],mul_res1[11519]);
multi_7x28 multi_7x28_mod_11520(clk,rst,matrix_A[11520],matrix_B[120],mul_res1[11520]);
multi_7x28 multi_7x28_mod_11521(clk,rst,matrix_A[11521],matrix_B[121],mul_res1[11521]);
multi_7x28 multi_7x28_mod_11522(clk,rst,matrix_A[11522],matrix_B[122],mul_res1[11522]);
multi_7x28 multi_7x28_mod_11523(clk,rst,matrix_A[11523],matrix_B[123],mul_res1[11523]);
multi_7x28 multi_7x28_mod_11524(clk,rst,matrix_A[11524],matrix_B[124],mul_res1[11524]);
multi_7x28 multi_7x28_mod_11525(clk,rst,matrix_A[11525],matrix_B[125],mul_res1[11525]);
multi_7x28 multi_7x28_mod_11526(clk,rst,matrix_A[11526],matrix_B[126],mul_res1[11526]);
multi_7x28 multi_7x28_mod_11527(clk,rst,matrix_A[11527],matrix_B[127],mul_res1[11527]);
multi_7x28 multi_7x28_mod_11528(clk,rst,matrix_A[11528],matrix_B[128],mul_res1[11528]);
multi_7x28 multi_7x28_mod_11529(clk,rst,matrix_A[11529],matrix_B[129],mul_res1[11529]);
multi_7x28 multi_7x28_mod_11530(clk,rst,matrix_A[11530],matrix_B[130],mul_res1[11530]);
multi_7x28 multi_7x28_mod_11531(clk,rst,matrix_A[11531],matrix_B[131],mul_res1[11531]);
multi_7x28 multi_7x28_mod_11532(clk,rst,matrix_A[11532],matrix_B[132],mul_res1[11532]);
multi_7x28 multi_7x28_mod_11533(clk,rst,matrix_A[11533],matrix_B[133],mul_res1[11533]);
multi_7x28 multi_7x28_mod_11534(clk,rst,matrix_A[11534],matrix_B[134],mul_res1[11534]);
multi_7x28 multi_7x28_mod_11535(clk,rst,matrix_A[11535],matrix_B[135],mul_res1[11535]);
multi_7x28 multi_7x28_mod_11536(clk,rst,matrix_A[11536],matrix_B[136],mul_res1[11536]);
multi_7x28 multi_7x28_mod_11537(clk,rst,matrix_A[11537],matrix_B[137],mul_res1[11537]);
multi_7x28 multi_7x28_mod_11538(clk,rst,matrix_A[11538],matrix_B[138],mul_res1[11538]);
multi_7x28 multi_7x28_mod_11539(clk,rst,matrix_A[11539],matrix_B[139],mul_res1[11539]);
multi_7x28 multi_7x28_mod_11540(clk,rst,matrix_A[11540],matrix_B[140],mul_res1[11540]);
multi_7x28 multi_7x28_mod_11541(clk,rst,matrix_A[11541],matrix_B[141],mul_res1[11541]);
multi_7x28 multi_7x28_mod_11542(clk,rst,matrix_A[11542],matrix_B[142],mul_res1[11542]);
multi_7x28 multi_7x28_mod_11543(clk,rst,matrix_A[11543],matrix_B[143],mul_res1[11543]);
multi_7x28 multi_7x28_mod_11544(clk,rst,matrix_A[11544],matrix_B[144],mul_res1[11544]);
multi_7x28 multi_7x28_mod_11545(clk,rst,matrix_A[11545],matrix_B[145],mul_res1[11545]);
multi_7x28 multi_7x28_mod_11546(clk,rst,matrix_A[11546],matrix_B[146],mul_res1[11546]);
multi_7x28 multi_7x28_mod_11547(clk,rst,matrix_A[11547],matrix_B[147],mul_res1[11547]);
multi_7x28 multi_7x28_mod_11548(clk,rst,matrix_A[11548],matrix_B[148],mul_res1[11548]);
multi_7x28 multi_7x28_mod_11549(clk,rst,matrix_A[11549],matrix_B[149],mul_res1[11549]);
multi_7x28 multi_7x28_mod_11550(clk,rst,matrix_A[11550],matrix_B[150],mul_res1[11550]);
multi_7x28 multi_7x28_mod_11551(clk,rst,matrix_A[11551],matrix_B[151],mul_res1[11551]);
multi_7x28 multi_7x28_mod_11552(clk,rst,matrix_A[11552],matrix_B[152],mul_res1[11552]);
multi_7x28 multi_7x28_mod_11553(clk,rst,matrix_A[11553],matrix_B[153],mul_res1[11553]);
multi_7x28 multi_7x28_mod_11554(clk,rst,matrix_A[11554],matrix_B[154],mul_res1[11554]);
multi_7x28 multi_7x28_mod_11555(clk,rst,matrix_A[11555],matrix_B[155],mul_res1[11555]);
multi_7x28 multi_7x28_mod_11556(clk,rst,matrix_A[11556],matrix_B[156],mul_res1[11556]);
multi_7x28 multi_7x28_mod_11557(clk,rst,matrix_A[11557],matrix_B[157],mul_res1[11557]);
multi_7x28 multi_7x28_mod_11558(clk,rst,matrix_A[11558],matrix_B[158],mul_res1[11558]);
multi_7x28 multi_7x28_mod_11559(clk,rst,matrix_A[11559],matrix_B[159],mul_res1[11559]);
multi_7x28 multi_7x28_mod_11560(clk,rst,matrix_A[11560],matrix_B[160],mul_res1[11560]);
multi_7x28 multi_7x28_mod_11561(clk,rst,matrix_A[11561],matrix_B[161],mul_res1[11561]);
multi_7x28 multi_7x28_mod_11562(clk,rst,matrix_A[11562],matrix_B[162],mul_res1[11562]);
multi_7x28 multi_7x28_mod_11563(clk,rst,matrix_A[11563],matrix_B[163],mul_res1[11563]);
multi_7x28 multi_7x28_mod_11564(clk,rst,matrix_A[11564],matrix_B[164],mul_res1[11564]);
multi_7x28 multi_7x28_mod_11565(clk,rst,matrix_A[11565],matrix_B[165],mul_res1[11565]);
multi_7x28 multi_7x28_mod_11566(clk,rst,matrix_A[11566],matrix_B[166],mul_res1[11566]);
multi_7x28 multi_7x28_mod_11567(clk,rst,matrix_A[11567],matrix_B[167],mul_res1[11567]);
multi_7x28 multi_7x28_mod_11568(clk,rst,matrix_A[11568],matrix_B[168],mul_res1[11568]);
multi_7x28 multi_7x28_mod_11569(clk,rst,matrix_A[11569],matrix_B[169],mul_res1[11569]);
multi_7x28 multi_7x28_mod_11570(clk,rst,matrix_A[11570],matrix_B[170],mul_res1[11570]);
multi_7x28 multi_7x28_mod_11571(clk,rst,matrix_A[11571],matrix_B[171],mul_res1[11571]);
multi_7x28 multi_7x28_mod_11572(clk,rst,matrix_A[11572],matrix_B[172],mul_res1[11572]);
multi_7x28 multi_7x28_mod_11573(clk,rst,matrix_A[11573],matrix_B[173],mul_res1[11573]);
multi_7x28 multi_7x28_mod_11574(clk,rst,matrix_A[11574],matrix_B[174],mul_res1[11574]);
multi_7x28 multi_7x28_mod_11575(clk,rst,matrix_A[11575],matrix_B[175],mul_res1[11575]);
multi_7x28 multi_7x28_mod_11576(clk,rst,matrix_A[11576],matrix_B[176],mul_res1[11576]);
multi_7x28 multi_7x28_mod_11577(clk,rst,matrix_A[11577],matrix_B[177],mul_res1[11577]);
multi_7x28 multi_7x28_mod_11578(clk,rst,matrix_A[11578],matrix_B[178],mul_res1[11578]);
multi_7x28 multi_7x28_mod_11579(clk,rst,matrix_A[11579],matrix_B[179],mul_res1[11579]);
multi_7x28 multi_7x28_mod_11580(clk,rst,matrix_A[11580],matrix_B[180],mul_res1[11580]);
multi_7x28 multi_7x28_mod_11581(clk,rst,matrix_A[11581],matrix_B[181],mul_res1[11581]);
multi_7x28 multi_7x28_mod_11582(clk,rst,matrix_A[11582],matrix_B[182],mul_res1[11582]);
multi_7x28 multi_7x28_mod_11583(clk,rst,matrix_A[11583],matrix_B[183],mul_res1[11583]);
multi_7x28 multi_7x28_mod_11584(clk,rst,matrix_A[11584],matrix_B[184],mul_res1[11584]);
multi_7x28 multi_7x28_mod_11585(clk,rst,matrix_A[11585],matrix_B[185],mul_res1[11585]);
multi_7x28 multi_7x28_mod_11586(clk,rst,matrix_A[11586],matrix_B[186],mul_res1[11586]);
multi_7x28 multi_7x28_mod_11587(clk,rst,matrix_A[11587],matrix_B[187],mul_res1[11587]);
multi_7x28 multi_7x28_mod_11588(clk,rst,matrix_A[11588],matrix_B[188],mul_res1[11588]);
multi_7x28 multi_7x28_mod_11589(clk,rst,matrix_A[11589],matrix_B[189],mul_res1[11589]);
multi_7x28 multi_7x28_mod_11590(clk,rst,matrix_A[11590],matrix_B[190],mul_res1[11590]);
multi_7x28 multi_7x28_mod_11591(clk,rst,matrix_A[11591],matrix_B[191],mul_res1[11591]);
multi_7x28 multi_7x28_mod_11592(clk,rst,matrix_A[11592],matrix_B[192],mul_res1[11592]);
multi_7x28 multi_7x28_mod_11593(clk,rst,matrix_A[11593],matrix_B[193],mul_res1[11593]);
multi_7x28 multi_7x28_mod_11594(clk,rst,matrix_A[11594],matrix_B[194],mul_res1[11594]);
multi_7x28 multi_7x28_mod_11595(clk,rst,matrix_A[11595],matrix_B[195],mul_res1[11595]);
multi_7x28 multi_7x28_mod_11596(clk,rst,matrix_A[11596],matrix_B[196],mul_res1[11596]);
multi_7x28 multi_7x28_mod_11597(clk,rst,matrix_A[11597],matrix_B[197],mul_res1[11597]);
multi_7x28 multi_7x28_mod_11598(clk,rst,matrix_A[11598],matrix_B[198],mul_res1[11598]);
multi_7x28 multi_7x28_mod_11599(clk,rst,matrix_A[11599],matrix_B[199],mul_res1[11599]);
multi_7x28 multi_7x28_mod_11600(clk,rst,matrix_A[11600],matrix_B[0],mul_res1[11600]);
multi_7x28 multi_7x28_mod_11601(clk,rst,matrix_A[11601],matrix_B[1],mul_res1[11601]);
multi_7x28 multi_7x28_mod_11602(clk,rst,matrix_A[11602],matrix_B[2],mul_res1[11602]);
multi_7x28 multi_7x28_mod_11603(clk,rst,matrix_A[11603],matrix_B[3],mul_res1[11603]);
multi_7x28 multi_7x28_mod_11604(clk,rst,matrix_A[11604],matrix_B[4],mul_res1[11604]);
multi_7x28 multi_7x28_mod_11605(clk,rst,matrix_A[11605],matrix_B[5],mul_res1[11605]);
multi_7x28 multi_7x28_mod_11606(clk,rst,matrix_A[11606],matrix_B[6],mul_res1[11606]);
multi_7x28 multi_7x28_mod_11607(clk,rst,matrix_A[11607],matrix_B[7],mul_res1[11607]);
multi_7x28 multi_7x28_mod_11608(clk,rst,matrix_A[11608],matrix_B[8],mul_res1[11608]);
multi_7x28 multi_7x28_mod_11609(clk,rst,matrix_A[11609],matrix_B[9],mul_res1[11609]);
multi_7x28 multi_7x28_mod_11610(clk,rst,matrix_A[11610],matrix_B[10],mul_res1[11610]);
multi_7x28 multi_7x28_mod_11611(clk,rst,matrix_A[11611],matrix_B[11],mul_res1[11611]);
multi_7x28 multi_7x28_mod_11612(clk,rst,matrix_A[11612],matrix_B[12],mul_res1[11612]);
multi_7x28 multi_7x28_mod_11613(clk,rst,matrix_A[11613],matrix_B[13],mul_res1[11613]);
multi_7x28 multi_7x28_mod_11614(clk,rst,matrix_A[11614],matrix_B[14],mul_res1[11614]);
multi_7x28 multi_7x28_mod_11615(clk,rst,matrix_A[11615],matrix_B[15],mul_res1[11615]);
multi_7x28 multi_7x28_mod_11616(clk,rst,matrix_A[11616],matrix_B[16],mul_res1[11616]);
multi_7x28 multi_7x28_mod_11617(clk,rst,matrix_A[11617],matrix_B[17],mul_res1[11617]);
multi_7x28 multi_7x28_mod_11618(clk,rst,matrix_A[11618],matrix_B[18],mul_res1[11618]);
multi_7x28 multi_7x28_mod_11619(clk,rst,matrix_A[11619],matrix_B[19],mul_res1[11619]);
multi_7x28 multi_7x28_mod_11620(clk,rst,matrix_A[11620],matrix_B[20],mul_res1[11620]);
multi_7x28 multi_7x28_mod_11621(clk,rst,matrix_A[11621],matrix_B[21],mul_res1[11621]);
multi_7x28 multi_7x28_mod_11622(clk,rst,matrix_A[11622],matrix_B[22],mul_res1[11622]);
multi_7x28 multi_7x28_mod_11623(clk,rst,matrix_A[11623],matrix_B[23],mul_res1[11623]);
multi_7x28 multi_7x28_mod_11624(clk,rst,matrix_A[11624],matrix_B[24],mul_res1[11624]);
multi_7x28 multi_7x28_mod_11625(clk,rst,matrix_A[11625],matrix_B[25],mul_res1[11625]);
multi_7x28 multi_7x28_mod_11626(clk,rst,matrix_A[11626],matrix_B[26],mul_res1[11626]);
multi_7x28 multi_7x28_mod_11627(clk,rst,matrix_A[11627],matrix_B[27],mul_res1[11627]);
multi_7x28 multi_7x28_mod_11628(clk,rst,matrix_A[11628],matrix_B[28],mul_res1[11628]);
multi_7x28 multi_7x28_mod_11629(clk,rst,matrix_A[11629],matrix_B[29],mul_res1[11629]);
multi_7x28 multi_7x28_mod_11630(clk,rst,matrix_A[11630],matrix_B[30],mul_res1[11630]);
multi_7x28 multi_7x28_mod_11631(clk,rst,matrix_A[11631],matrix_B[31],mul_res1[11631]);
multi_7x28 multi_7x28_mod_11632(clk,rst,matrix_A[11632],matrix_B[32],mul_res1[11632]);
multi_7x28 multi_7x28_mod_11633(clk,rst,matrix_A[11633],matrix_B[33],mul_res1[11633]);
multi_7x28 multi_7x28_mod_11634(clk,rst,matrix_A[11634],matrix_B[34],mul_res1[11634]);
multi_7x28 multi_7x28_mod_11635(clk,rst,matrix_A[11635],matrix_B[35],mul_res1[11635]);
multi_7x28 multi_7x28_mod_11636(clk,rst,matrix_A[11636],matrix_B[36],mul_res1[11636]);
multi_7x28 multi_7x28_mod_11637(clk,rst,matrix_A[11637],matrix_B[37],mul_res1[11637]);
multi_7x28 multi_7x28_mod_11638(clk,rst,matrix_A[11638],matrix_B[38],mul_res1[11638]);
multi_7x28 multi_7x28_mod_11639(clk,rst,matrix_A[11639],matrix_B[39],mul_res1[11639]);
multi_7x28 multi_7x28_mod_11640(clk,rst,matrix_A[11640],matrix_B[40],mul_res1[11640]);
multi_7x28 multi_7x28_mod_11641(clk,rst,matrix_A[11641],matrix_B[41],mul_res1[11641]);
multi_7x28 multi_7x28_mod_11642(clk,rst,matrix_A[11642],matrix_B[42],mul_res1[11642]);
multi_7x28 multi_7x28_mod_11643(clk,rst,matrix_A[11643],matrix_B[43],mul_res1[11643]);
multi_7x28 multi_7x28_mod_11644(clk,rst,matrix_A[11644],matrix_B[44],mul_res1[11644]);
multi_7x28 multi_7x28_mod_11645(clk,rst,matrix_A[11645],matrix_B[45],mul_res1[11645]);
multi_7x28 multi_7x28_mod_11646(clk,rst,matrix_A[11646],matrix_B[46],mul_res1[11646]);
multi_7x28 multi_7x28_mod_11647(clk,rst,matrix_A[11647],matrix_B[47],mul_res1[11647]);
multi_7x28 multi_7x28_mod_11648(clk,rst,matrix_A[11648],matrix_B[48],mul_res1[11648]);
multi_7x28 multi_7x28_mod_11649(clk,rst,matrix_A[11649],matrix_B[49],mul_res1[11649]);
multi_7x28 multi_7x28_mod_11650(clk,rst,matrix_A[11650],matrix_B[50],mul_res1[11650]);
multi_7x28 multi_7x28_mod_11651(clk,rst,matrix_A[11651],matrix_B[51],mul_res1[11651]);
multi_7x28 multi_7x28_mod_11652(clk,rst,matrix_A[11652],matrix_B[52],mul_res1[11652]);
multi_7x28 multi_7x28_mod_11653(clk,rst,matrix_A[11653],matrix_B[53],mul_res1[11653]);
multi_7x28 multi_7x28_mod_11654(clk,rst,matrix_A[11654],matrix_B[54],mul_res1[11654]);
multi_7x28 multi_7x28_mod_11655(clk,rst,matrix_A[11655],matrix_B[55],mul_res1[11655]);
multi_7x28 multi_7x28_mod_11656(clk,rst,matrix_A[11656],matrix_B[56],mul_res1[11656]);
multi_7x28 multi_7x28_mod_11657(clk,rst,matrix_A[11657],matrix_B[57],mul_res1[11657]);
multi_7x28 multi_7x28_mod_11658(clk,rst,matrix_A[11658],matrix_B[58],mul_res1[11658]);
multi_7x28 multi_7x28_mod_11659(clk,rst,matrix_A[11659],matrix_B[59],mul_res1[11659]);
multi_7x28 multi_7x28_mod_11660(clk,rst,matrix_A[11660],matrix_B[60],mul_res1[11660]);
multi_7x28 multi_7x28_mod_11661(clk,rst,matrix_A[11661],matrix_B[61],mul_res1[11661]);
multi_7x28 multi_7x28_mod_11662(clk,rst,matrix_A[11662],matrix_B[62],mul_res1[11662]);
multi_7x28 multi_7x28_mod_11663(clk,rst,matrix_A[11663],matrix_B[63],mul_res1[11663]);
multi_7x28 multi_7x28_mod_11664(clk,rst,matrix_A[11664],matrix_B[64],mul_res1[11664]);
multi_7x28 multi_7x28_mod_11665(clk,rst,matrix_A[11665],matrix_B[65],mul_res1[11665]);
multi_7x28 multi_7x28_mod_11666(clk,rst,matrix_A[11666],matrix_B[66],mul_res1[11666]);
multi_7x28 multi_7x28_mod_11667(clk,rst,matrix_A[11667],matrix_B[67],mul_res1[11667]);
multi_7x28 multi_7x28_mod_11668(clk,rst,matrix_A[11668],matrix_B[68],mul_res1[11668]);
multi_7x28 multi_7x28_mod_11669(clk,rst,matrix_A[11669],matrix_B[69],mul_res1[11669]);
multi_7x28 multi_7x28_mod_11670(clk,rst,matrix_A[11670],matrix_B[70],mul_res1[11670]);
multi_7x28 multi_7x28_mod_11671(clk,rst,matrix_A[11671],matrix_B[71],mul_res1[11671]);
multi_7x28 multi_7x28_mod_11672(clk,rst,matrix_A[11672],matrix_B[72],mul_res1[11672]);
multi_7x28 multi_7x28_mod_11673(clk,rst,matrix_A[11673],matrix_B[73],mul_res1[11673]);
multi_7x28 multi_7x28_mod_11674(clk,rst,matrix_A[11674],matrix_B[74],mul_res1[11674]);
multi_7x28 multi_7x28_mod_11675(clk,rst,matrix_A[11675],matrix_B[75],mul_res1[11675]);
multi_7x28 multi_7x28_mod_11676(clk,rst,matrix_A[11676],matrix_B[76],mul_res1[11676]);
multi_7x28 multi_7x28_mod_11677(clk,rst,matrix_A[11677],matrix_B[77],mul_res1[11677]);
multi_7x28 multi_7x28_mod_11678(clk,rst,matrix_A[11678],matrix_B[78],mul_res1[11678]);
multi_7x28 multi_7x28_mod_11679(clk,rst,matrix_A[11679],matrix_B[79],mul_res1[11679]);
multi_7x28 multi_7x28_mod_11680(clk,rst,matrix_A[11680],matrix_B[80],mul_res1[11680]);
multi_7x28 multi_7x28_mod_11681(clk,rst,matrix_A[11681],matrix_B[81],mul_res1[11681]);
multi_7x28 multi_7x28_mod_11682(clk,rst,matrix_A[11682],matrix_B[82],mul_res1[11682]);
multi_7x28 multi_7x28_mod_11683(clk,rst,matrix_A[11683],matrix_B[83],mul_res1[11683]);
multi_7x28 multi_7x28_mod_11684(clk,rst,matrix_A[11684],matrix_B[84],mul_res1[11684]);
multi_7x28 multi_7x28_mod_11685(clk,rst,matrix_A[11685],matrix_B[85],mul_res1[11685]);
multi_7x28 multi_7x28_mod_11686(clk,rst,matrix_A[11686],matrix_B[86],mul_res1[11686]);
multi_7x28 multi_7x28_mod_11687(clk,rst,matrix_A[11687],matrix_B[87],mul_res1[11687]);
multi_7x28 multi_7x28_mod_11688(clk,rst,matrix_A[11688],matrix_B[88],mul_res1[11688]);
multi_7x28 multi_7x28_mod_11689(clk,rst,matrix_A[11689],matrix_B[89],mul_res1[11689]);
multi_7x28 multi_7x28_mod_11690(clk,rst,matrix_A[11690],matrix_B[90],mul_res1[11690]);
multi_7x28 multi_7x28_mod_11691(clk,rst,matrix_A[11691],matrix_B[91],mul_res1[11691]);
multi_7x28 multi_7x28_mod_11692(clk,rst,matrix_A[11692],matrix_B[92],mul_res1[11692]);
multi_7x28 multi_7x28_mod_11693(clk,rst,matrix_A[11693],matrix_B[93],mul_res1[11693]);
multi_7x28 multi_7x28_mod_11694(clk,rst,matrix_A[11694],matrix_B[94],mul_res1[11694]);
multi_7x28 multi_7x28_mod_11695(clk,rst,matrix_A[11695],matrix_B[95],mul_res1[11695]);
multi_7x28 multi_7x28_mod_11696(clk,rst,matrix_A[11696],matrix_B[96],mul_res1[11696]);
multi_7x28 multi_7x28_mod_11697(clk,rst,matrix_A[11697],matrix_B[97],mul_res1[11697]);
multi_7x28 multi_7x28_mod_11698(clk,rst,matrix_A[11698],matrix_B[98],mul_res1[11698]);
multi_7x28 multi_7x28_mod_11699(clk,rst,matrix_A[11699],matrix_B[99],mul_res1[11699]);
multi_7x28 multi_7x28_mod_11700(clk,rst,matrix_A[11700],matrix_B[100],mul_res1[11700]);
multi_7x28 multi_7x28_mod_11701(clk,rst,matrix_A[11701],matrix_B[101],mul_res1[11701]);
multi_7x28 multi_7x28_mod_11702(clk,rst,matrix_A[11702],matrix_B[102],mul_res1[11702]);
multi_7x28 multi_7x28_mod_11703(clk,rst,matrix_A[11703],matrix_B[103],mul_res1[11703]);
multi_7x28 multi_7x28_mod_11704(clk,rst,matrix_A[11704],matrix_B[104],mul_res1[11704]);
multi_7x28 multi_7x28_mod_11705(clk,rst,matrix_A[11705],matrix_B[105],mul_res1[11705]);
multi_7x28 multi_7x28_mod_11706(clk,rst,matrix_A[11706],matrix_B[106],mul_res1[11706]);
multi_7x28 multi_7x28_mod_11707(clk,rst,matrix_A[11707],matrix_B[107],mul_res1[11707]);
multi_7x28 multi_7x28_mod_11708(clk,rst,matrix_A[11708],matrix_B[108],mul_res1[11708]);
multi_7x28 multi_7x28_mod_11709(clk,rst,matrix_A[11709],matrix_B[109],mul_res1[11709]);
multi_7x28 multi_7x28_mod_11710(clk,rst,matrix_A[11710],matrix_B[110],mul_res1[11710]);
multi_7x28 multi_7x28_mod_11711(clk,rst,matrix_A[11711],matrix_B[111],mul_res1[11711]);
multi_7x28 multi_7x28_mod_11712(clk,rst,matrix_A[11712],matrix_B[112],mul_res1[11712]);
multi_7x28 multi_7x28_mod_11713(clk,rst,matrix_A[11713],matrix_B[113],mul_res1[11713]);
multi_7x28 multi_7x28_mod_11714(clk,rst,matrix_A[11714],matrix_B[114],mul_res1[11714]);
multi_7x28 multi_7x28_mod_11715(clk,rst,matrix_A[11715],matrix_B[115],mul_res1[11715]);
multi_7x28 multi_7x28_mod_11716(clk,rst,matrix_A[11716],matrix_B[116],mul_res1[11716]);
multi_7x28 multi_7x28_mod_11717(clk,rst,matrix_A[11717],matrix_B[117],mul_res1[11717]);
multi_7x28 multi_7x28_mod_11718(clk,rst,matrix_A[11718],matrix_B[118],mul_res1[11718]);
multi_7x28 multi_7x28_mod_11719(clk,rst,matrix_A[11719],matrix_B[119],mul_res1[11719]);
multi_7x28 multi_7x28_mod_11720(clk,rst,matrix_A[11720],matrix_B[120],mul_res1[11720]);
multi_7x28 multi_7x28_mod_11721(clk,rst,matrix_A[11721],matrix_B[121],mul_res1[11721]);
multi_7x28 multi_7x28_mod_11722(clk,rst,matrix_A[11722],matrix_B[122],mul_res1[11722]);
multi_7x28 multi_7x28_mod_11723(clk,rst,matrix_A[11723],matrix_B[123],mul_res1[11723]);
multi_7x28 multi_7x28_mod_11724(clk,rst,matrix_A[11724],matrix_B[124],mul_res1[11724]);
multi_7x28 multi_7x28_mod_11725(clk,rst,matrix_A[11725],matrix_B[125],mul_res1[11725]);
multi_7x28 multi_7x28_mod_11726(clk,rst,matrix_A[11726],matrix_B[126],mul_res1[11726]);
multi_7x28 multi_7x28_mod_11727(clk,rst,matrix_A[11727],matrix_B[127],mul_res1[11727]);
multi_7x28 multi_7x28_mod_11728(clk,rst,matrix_A[11728],matrix_B[128],mul_res1[11728]);
multi_7x28 multi_7x28_mod_11729(clk,rst,matrix_A[11729],matrix_B[129],mul_res1[11729]);
multi_7x28 multi_7x28_mod_11730(clk,rst,matrix_A[11730],matrix_B[130],mul_res1[11730]);
multi_7x28 multi_7x28_mod_11731(clk,rst,matrix_A[11731],matrix_B[131],mul_res1[11731]);
multi_7x28 multi_7x28_mod_11732(clk,rst,matrix_A[11732],matrix_B[132],mul_res1[11732]);
multi_7x28 multi_7x28_mod_11733(clk,rst,matrix_A[11733],matrix_B[133],mul_res1[11733]);
multi_7x28 multi_7x28_mod_11734(clk,rst,matrix_A[11734],matrix_B[134],mul_res1[11734]);
multi_7x28 multi_7x28_mod_11735(clk,rst,matrix_A[11735],matrix_B[135],mul_res1[11735]);
multi_7x28 multi_7x28_mod_11736(clk,rst,matrix_A[11736],matrix_B[136],mul_res1[11736]);
multi_7x28 multi_7x28_mod_11737(clk,rst,matrix_A[11737],matrix_B[137],mul_res1[11737]);
multi_7x28 multi_7x28_mod_11738(clk,rst,matrix_A[11738],matrix_B[138],mul_res1[11738]);
multi_7x28 multi_7x28_mod_11739(clk,rst,matrix_A[11739],matrix_B[139],mul_res1[11739]);
multi_7x28 multi_7x28_mod_11740(clk,rst,matrix_A[11740],matrix_B[140],mul_res1[11740]);
multi_7x28 multi_7x28_mod_11741(clk,rst,matrix_A[11741],matrix_B[141],mul_res1[11741]);
multi_7x28 multi_7x28_mod_11742(clk,rst,matrix_A[11742],matrix_B[142],mul_res1[11742]);
multi_7x28 multi_7x28_mod_11743(clk,rst,matrix_A[11743],matrix_B[143],mul_res1[11743]);
multi_7x28 multi_7x28_mod_11744(clk,rst,matrix_A[11744],matrix_B[144],mul_res1[11744]);
multi_7x28 multi_7x28_mod_11745(clk,rst,matrix_A[11745],matrix_B[145],mul_res1[11745]);
multi_7x28 multi_7x28_mod_11746(clk,rst,matrix_A[11746],matrix_B[146],mul_res1[11746]);
multi_7x28 multi_7x28_mod_11747(clk,rst,matrix_A[11747],matrix_B[147],mul_res1[11747]);
multi_7x28 multi_7x28_mod_11748(clk,rst,matrix_A[11748],matrix_B[148],mul_res1[11748]);
multi_7x28 multi_7x28_mod_11749(clk,rst,matrix_A[11749],matrix_B[149],mul_res1[11749]);
multi_7x28 multi_7x28_mod_11750(clk,rst,matrix_A[11750],matrix_B[150],mul_res1[11750]);
multi_7x28 multi_7x28_mod_11751(clk,rst,matrix_A[11751],matrix_B[151],mul_res1[11751]);
multi_7x28 multi_7x28_mod_11752(clk,rst,matrix_A[11752],matrix_B[152],mul_res1[11752]);
multi_7x28 multi_7x28_mod_11753(clk,rst,matrix_A[11753],matrix_B[153],mul_res1[11753]);
multi_7x28 multi_7x28_mod_11754(clk,rst,matrix_A[11754],matrix_B[154],mul_res1[11754]);
multi_7x28 multi_7x28_mod_11755(clk,rst,matrix_A[11755],matrix_B[155],mul_res1[11755]);
multi_7x28 multi_7x28_mod_11756(clk,rst,matrix_A[11756],matrix_B[156],mul_res1[11756]);
multi_7x28 multi_7x28_mod_11757(clk,rst,matrix_A[11757],matrix_B[157],mul_res1[11757]);
multi_7x28 multi_7x28_mod_11758(clk,rst,matrix_A[11758],matrix_B[158],mul_res1[11758]);
multi_7x28 multi_7x28_mod_11759(clk,rst,matrix_A[11759],matrix_B[159],mul_res1[11759]);
multi_7x28 multi_7x28_mod_11760(clk,rst,matrix_A[11760],matrix_B[160],mul_res1[11760]);
multi_7x28 multi_7x28_mod_11761(clk,rst,matrix_A[11761],matrix_B[161],mul_res1[11761]);
multi_7x28 multi_7x28_mod_11762(clk,rst,matrix_A[11762],matrix_B[162],mul_res1[11762]);
multi_7x28 multi_7x28_mod_11763(clk,rst,matrix_A[11763],matrix_B[163],mul_res1[11763]);
multi_7x28 multi_7x28_mod_11764(clk,rst,matrix_A[11764],matrix_B[164],mul_res1[11764]);
multi_7x28 multi_7x28_mod_11765(clk,rst,matrix_A[11765],matrix_B[165],mul_res1[11765]);
multi_7x28 multi_7x28_mod_11766(clk,rst,matrix_A[11766],matrix_B[166],mul_res1[11766]);
multi_7x28 multi_7x28_mod_11767(clk,rst,matrix_A[11767],matrix_B[167],mul_res1[11767]);
multi_7x28 multi_7x28_mod_11768(clk,rst,matrix_A[11768],matrix_B[168],mul_res1[11768]);
multi_7x28 multi_7x28_mod_11769(clk,rst,matrix_A[11769],matrix_B[169],mul_res1[11769]);
multi_7x28 multi_7x28_mod_11770(clk,rst,matrix_A[11770],matrix_B[170],mul_res1[11770]);
multi_7x28 multi_7x28_mod_11771(clk,rst,matrix_A[11771],matrix_B[171],mul_res1[11771]);
multi_7x28 multi_7x28_mod_11772(clk,rst,matrix_A[11772],matrix_B[172],mul_res1[11772]);
multi_7x28 multi_7x28_mod_11773(clk,rst,matrix_A[11773],matrix_B[173],mul_res1[11773]);
multi_7x28 multi_7x28_mod_11774(clk,rst,matrix_A[11774],matrix_B[174],mul_res1[11774]);
multi_7x28 multi_7x28_mod_11775(clk,rst,matrix_A[11775],matrix_B[175],mul_res1[11775]);
multi_7x28 multi_7x28_mod_11776(clk,rst,matrix_A[11776],matrix_B[176],mul_res1[11776]);
multi_7x28 multi_7x28_mod_11777(clk,rst,matrix_A[11777],matrix_B[177],mul_res1[11777]);
multi_7x28 multi_7x28_mod_11778(clk,rst,matrix_A[11778],matrix_B[178],mul_res1[11778]);
multi_7x28 multi_7x28_mod_11779(clk,rst,matrix_A[11779],matrix_B[179],mul_res1[11779]);
multi_7x28 multi_7x28_mod_11780(clk,rst,matrix_A[11780],matrix_B[180],mul_res1[11780]);
multi_7x28 multi_7x28_mod_11781(clk,rst,matrix_A[11781],matrix_B[181],mul_res1[11781]);
multi_7x28 multi_7x28_mod_11782(clk,rst,matrix_A[11782],matrix_B[182],mul_res1[11782]);
multi_7x28 multi_7x28_mod_11783(clk,rst,matrix_A[11783],matrix_B[183],mul_res1[11783]);
multi_7x28 multi_7x28_mod_11784(clk,rst,matrix_A[11784],matrix_B[184],mul_res1[11784]);
multi_7x28 multi_7x28_mod_11785(clk,rst,matrix_A[11785],matrix_B[185],mul_res1[11785]);
multi_7x28 multi_7x28_mod_11786(clk,rst,matrix_A[11786],matrix_B[186],mul_res1[11786]);
multi_7x28 multi_7x28_mod_11787(clk,rst,matrix_A[11787],matrix_B[187],mul_res1[11787]);
multi_7x28 multi_7x28_mod_11788(clk,rst,matrix_A[11788],matrix_B[188],mul_res1[11788]);
multi_7x28 multi_7x28_mod_11789(clk,rst,matrix_A[11789],matrix_B[189],mul_res1[11789]);
multi_7x28 multi_7x28_mod_11790(clk,rst,matrix_A[11790],matrix_B[190],mul_res1[11790]);
multi_7x28 multi_7x28_mod_11791(clk,rst,matrix_A[11791],matrix_B[191],mul_res1[11791]);
multi_7x28 multi_7x28_mod_11792(clk,rst,matrix_A[11792],matrix_B[192],mul_res1[11792]);
multi_7x28 multi_7x28_mod_11793(clk,rst,matrix_A[11793],matrix_B[193],mul_res1[11793]);
multi_7x28 multi_7x28_mod_11794(clk,rst,matrix_A[11794],matrix_B[194],mul_res1[11794]);
multi_7x28 multi_7x28_mod_11795(clk,rst,matrix_A[11795],matrix_B[195],mul_res1[11795]);
multi_7x28 multi_7x28_mod_11796(clk,rst,matrix_A[11796],matrix_B[196],mul_res1[11796]);
multi_7x28 multi_7x28_mod_11797(clk,rst,matrix_A[11797],matrix_B[197],mul_res1[11797]);
multi_7x28 multi_7x28_mod_11798(clk,rst,matrix_A[11798],matrix_B[198],mul_res1[11798]);
multi_7x28 multi_7x28_mod_11799(clk,rst,matrix_A[11799],matrix_B[199],mul_res1[11799]);
multi_7x28 multi_7x28_mod_11800(clk,rst,matrix_A[11800],matrix_B[0],mul_res1[11800]);
multi_7x28 multi_7x28_mod_11801(clk,rst,matrix_A[11801],matrix_B[1],mul_res1[11801]);
multi_7x28 multi_7x28_mod_11802(clk,rst,matrix_A[11802],matrix_B[2],mul_res1[11802]);
multi_7x28 multi_7x28_mod_11803(clk,rst,matrix_A[11803],matrix_B[3],mul_res1[11803]);
multi_7x28 multi_7x28_mod_11804(clk,rst,matrix_A[11804],matrix_B[4],mul_res1[11804]);
multi_7x28 multi_7x28_mod_11805(clk,rst,matrix_A[11805],matrix_B[5],mul_res1[11805]);
multi_7x28 multi_7x28_mod_11806(clk,rst,matrix_A[11806],matrix_B[6],mul_res1[11806]);
multi_7x28 multi_7x28_mod_11807(clk,rst,matrix_A[11807],matrix_B[7],mul_res1[11807]);
multi_7x28 multi_7x28_mod_11808(clk,rst,matrix_A[11808],matrix_B[8],mul_res1[11808]);
multi_7x28 multi_7x28_mod_11809(clk,rst,matrix_A[11809],matrix_B[9],mul_res1[11809]);
multi_7x28 multi_7x28_mod_11810(clk,rst,matrix_A[11810],matrix_B[10],mul_res1[11810]);
multi_7x28 multi_7x28_mod_11811(clk,rst,matrix_A[11811],matrix_B[11],mul_res1[11811]);
multi_7x28 multi_7x28_mod_11812(clk,rst,matrix_A[11812],matrix_B[12],mul_res1[11812]);
multi_7x28 multi_7x28_mod_11813(clk,rst,matrix_A[11813],matrix_B[13],mul_res1[11813]);
multi_7x28 multi_7x28_mod_11814(clk,rst,matrix_A[11814],matrix_B[14],mul_res1[11814]);
multi_7x28 multi_7x28_mod_11815(clk,rst,matrix_A[11815],matrix_B[15],mul_res1[11815]);
multi_7x28 multi_7x28_mod_11816(clk,rst,matrix_A[11816],matrix_B[16],mul_res1[11816]);
multi_7x28 multi_7x28_mod_11817(clk,rst,matrix_A[11817],matrix_B[17],mul_res1[11817]);
multi_7x28 multi_7x28_mod_11818(clk,rst,matrix_A[11818],matrix_B[18],mul_res1[11818]);
multi_7x28 multi_7x28_mod_11819(clk,rst,matrix_A[11819],matrix_B[19],mul_res1[11819]);
multi_7x28 multi_7x28_mod_11820(clk,rst,matrix_A[11820],matrix_B[20],mul_res1[11820]);
multi_7x28 multi_7x28_mod_11821(clk,rst,matrix_A[11821],matrix_B[21],mul_res1[11821]);
multi_7x28 multi_7x28_mod_11822(clk,rst,matrix_A[11822],matrix_B[22],mul_res1[11822]);
multi_7x28 multi_7x28_mod_11823(clk,rst,matrix_A[11823],matrix_B[23],mul_res1[11823]);
multi_7x28 multi_7x28_mod_11824(clk,rst,matrix_A[11824],matrix_B[24],mul_res1[11824]);
multi_7x28 multi_7x28_mod_11825(clk,rst,matrix_A[11825],matrix_B[25],mul_res1[11825]);
multi_7x28 multi_7x28_mod_11826(clk,rst,matrix_A[11826],matrix_B[26],mul_res1[11826]);
multi_7x28 multi_7x28_mod_11827(clk,rst,matrix_A[11827],matrix_B[27],mul_res1[11827]);
multi_7x28 multi_7x28_mod_11828(clk,rst,matrix_A[11828],matrix_B[28],mul_res1[11828]);
multi_7x28 multi_7x28_mod_11829(clk,rst,matrix_A[11829],matrix_B[29],mul_res1[11829]);
multi_7x28 multi_7x28_mod_11830(clk,rst,matrix_A[11830],matrix_B[30],mul_res1[11830]);
multi_7x28 multi_7x28_mod_11831(clk,rst,matrix_A[11831],matrix_B[31],mul_res1[11831]);
multi_7x28 multi_7x28_mod_11832(clk,rst,matrix_A[11832],matrix_B[32],mul_res1[11832]);
multi_7x28 multi_7x28_mod_11833(clk,rst,matrix_A[11833],matrix_B[33],mul_res1[11833]);
multi_7x28 multi_7x28_mod_11834(clk,rst,matrix_A[11834],matrix_B[34],mul_res1[11834]);
multi_7x28 multi_7x28_mod_11835(clk,rst,matrix_A[11835],matrix_B[35],mul_res1[11835]);
multi_7x28 multi_7x28_mod_11836(clk,rst,matrix_A[11836],matrix_B[36],mul_res1[11836]);
multi_7x28 multi_7x28_mod_11837(clk,rst,matrix_A[11837],matrix_B[37],mul_res1[11837]);
multi_7x28 multi_7x28_mod_11838(clk,rst,matrix_A[11838],matrix_B[38],mul_res1[11838]);
multi_7x28 multi_7x28_mod_11839(clk,rst,matrix_A[11839],matrix_B[39],mul_res1[11839]);
multi_7x28 multi_7x28_mod_11840(clk,rst,matrix_A[11840],matrix_B[40],mul_res1[11840]);
multi_7x28 multi_7x28_mod_11841(clk,rst,matrix_A[11841],matrix_B[41],mul_res1[11841]);
multi_7x28 multi_7x28_mod_11842(clk,rst,matrix_A[11842],matrix_B[42],mul_res1[11842]);
multi_7x28 multi_7x28_mod_11843(clk,rst,matrix_A[11843],matrix_B[43],mul_res1[11843]);
multi_7x28 multi_7x28_mod_11844(clk,rst,matrix_A[11844],matrix_B[44],mul_res1[11844]);
multi_7x28 multi_7x28_mod_11845(clk,rst,matrix_A[11845],matrix_B[45],mul_res1[11845]);
multi_7x28 multi_7x28_mod_11846(clk,rst,matrix_A[11846],matrix_B[46],mul_res1[11846]);
multi_7x28 multi_7x28_mod_11847(clk,rst,matrix_A[11847],matrix_B[47],mul_res1[11847]);
multi_7x28 multi_7x28_mod_11848(clk,rst,matrix_A[11848],matrix_B[48],mul_res1[11848]);
multi_7x28 multi_7x28_mod_11849(clk,rst,matrix_A[11849],matrix_B[49],mul_res1[11849]);
multi_7x28 multi_7x28_mod_11850(clk,rst,matrix_A[11850],matrix_B[50],mul_res1[11850]);
multi_7x28 multi_7x28_mod_11851(clk,rst,matrix_A[11851],matrix_B[51],mul_res1[11851]);
multi_7x28 multi_7x28_mod_11852(clk,rst,matrix_A[11852],matrix_B[52],mul_res1[11852]);
multi_7x28 multi_7x28_mod_11853(clk,rst,matrix_A[11853],matrix_B[53],mul_res1[11853]);
multi_7x28 multi_7x28_mod_11854(clk,rst,matrix_A[11854],matrix_B[54],mul_res1[11854]);
multi_7x28 multi_7x28_mod_11855(clk,rst,matrix_A[11855],matrix_B[55],mul_res1[11855]);
multi_7x28 multi_7x28_mod_11856(clk,rst,matrix_A[11856],matrix_B[56],mul_res1[11856]);
multi_7x28 multi_7x28_mod_11857(clk,rst,matrix_A[11857],matrix_B[57],mul_res1[11857]);
multi_7x28 multi_7x28_mod_11858(clk,rst,matrix_A[11858],matrix_B[58],mul_res1[11858]);
multi_7x28 multi_7x28_mod_11859(clk,rst,matrix_A[11859],matrix_B[59],mul_res1[11859]);
multi_7x28 multi_7x28_mod_11860(clk,rst,matrix_A[11860],matrix_B[60],mul_res1[11860]);
multi_7x28 multi_7x28_mod_11861(clk,rst,matrix_A[11861],matrix_B[61],mul_res1[11861]);
multi_7x28 multi_7x28_mod_11862(clk,rst,matrix_A[11862],matrix_B[62],mul_res1[11862]);
multi_7x28 multi_7x28_mod_11863(clk,rst,matrix_A[11863],matrix_B[63],mul_res1[11863]);
multi_7x28 multi_7x28_mod_11864(clk,rst,matrix_A[11864],matrix_B[64],mul_res1[11864]);
multi_7x28 multi_7x28_mod_11865(clk,rst,matrix_A[11865],matrix_B[65],mul_res1[11865]);
multi_7x28 multi_7x28_mod_11866(clk,rst,matrix_A[11866],matrix_B[66],mul_res1[11866]);
multi_7x28 multi_7x28_mod_11867(clk,rst,matrix_A[11867],matrix_B[67],mul_res1[11867]);
multi_7x28 multi_7x28_mod_11868(clk,rst,matrix_A[11868],matrix_B[68],mul_res1[11868]);
multi_7x28 multi_7x28_mod_11869(clk,rst,matrix_A[11869],matrix_B[69],mul_res1[11869]);
multi_7x28 multi_7x28_mod_11870(clk,rst,matrix_A[11870],matrix_B[70],mul_res1[11870]);
multi_7x28 multi_7x28_mod_11871(clk,rst,matrix_A[11871],matrix_B[71],mul_res1[11871]);
multi_7x28 multi_7x28_mod_11872(clk,rst,matrix_A[11872],matrix_B[72],mul_res1[11872]);
multi_7x28 multi_7x28_mod_11873(clk,rst,matrix_A[11873],matrix_B[73],mul_res1[11873]);
multi_7x28 multi_7x28_mod_11874(clk,rst,matrix_A[11874],matrix_B[74],mul_res1[11874]);
multi_7x28 multi_7x28_mod_11875(clk,rst,matrix_A[11875],matrix_B[75],mul_res1[11875]);
multi_7x28 multi_7x28_mod_11876(clk,rst,matrix_A[11876],matrix_B[76],mul_res1[11876]);
multi_7x28 multi_7x28_mod_11877(clk,rst,matrix_A[11877],matrix_B[77],mul_res1[11877]);
multi_7x28 multi_7x28_mod_11878(clk,rst,matrix_A[11878],matrix_B[78],mul_res1[11878]);
multi_7x28 multi_7x28_mod_11879(clk,rst,matrix_A[11879],matrix_B[79],mul_res1[11879]);
multi_7x28 multi_7x28_mod_11880(clk,rst,matrix_A[11880],matrix_B[80],mul_res1[11880]);
multi_7x28 multi_7x28_mod_11881(clk,rst,matrix_A[11881],matrix_B[81],mul_res1[11881]);
multi_7x28 multi_7x28_mod_11882(clk,rst,matrix_A[11882],matrix_B[82],mul_res1[11882]);
multi_7x28 multi_7x28_mod_11883(clk,rst,matrix_A[11883],matrix_B[83],mul_res1[11883]);
multi_7x28 multi_7x28_mod_11884(clk,rst,matrix_A[11884],matrix_B[84],mul_res1[11884]);
multi_7x28 multi_7x28_mod_11885(clk,rst,matrix_A[11885],matrix_B[85],mul_res1[11885]);
multi_7x28 multi_7x28_mod_11886(clk,rst,matrix_A[11886],matrix_B[86],mul_res1[11886]);
multi_7x28 multi_7x28_mod_11887(clk,rst,matrix_A[11887],matrix_B[87],mul_res1[11887]);
multi_7x28 multi_7x28_mod_11888(clk,rst,matrix_A[11888],matrix_B[88],mul_res1[11888]);
multi_7x28 multi_7x28_mod_11889(clk,rst,matrix_A[11889],matrix_B[89],mul_res1[11889]);
multi_7x28 multi_7x28_mod_11890(clk,rst,matrix_A[11890],matrix_B[90],mul_res1[11890]);
multi_7x28 multi_7x28_mod_11891(clk,rst,matrix_A[11891],matrix_B[91],mul_res1[11891]);
multi_7x28 multi_7x28_mod_11892(clk,rst,matrix_A[11892],matrix_B[92],mul_res1[11892]);
multi_7x28 multi_7x28_mod_11893(clk,rst,matrix_A[11893],matrix_B[93],mul_res1[11893]);
multi_7x28 multi_7x28_mod_11894(clk,rst,matrix_A[11894],matrix_B[94],mul_res1[11894]);
multi_7x28 multi_7x28_mod_11895(clk,rst,matrix_A[11895],matrix_B[95],mul_res1[11895]);
multi_7x28 multi_7x28_mod_11896(clk,rst,matrix_A[11896],matrix_B[96],mul_res1[11896]);
multi_7x28 multi_7x28_mod_11897(clk,rst,matrix_A[11897],matrix_B[97],mul_res1[11897]);
multi_7x28 multi_7x28_mod_11898(clk,rst,matrix_A[11898],matrix_B[98],mul_res1[11898]);
multi_7x28 multi_7x28_mod_11899(clk,rst,matrix_A[11899],matrix_B[99],mul_res1[11899]);
multi_7x28 multi_7x28_mod_11900(clk,rst,matrix_A[11900],matrix_B[100],mul_res1[11900]);
multi_7x28 multi_7x28_mod_11901(clk,rst,matrix_A[11901],matrix_B[101],mul_res1[11901]);
multi_7x28 multi_7x28_mod_11902(clk,rst,matrix_A[11902],matrix_B[102],mul_res1[11902]);
multi_7x28 multi_7x28_mod_11903(clk,rst,matrix_A[11903],matrix_B[103],mul_res1[11903]);
multi_7x28 multi_7x28_mod_11904(clk,rst,matrix_A[11904],matrix_B[104],mul_res1[11904]);
multi_7x28 multi_7x28_mod_11905(clk,rst,matrix_A[11905],matrix_B[105],mul_res1[11905]);
multi_7x28 multi_7x28_mod_11906(clk,rst,matrix_A[11906],matrix_B[106],mul_res1[11906]);
multi_7x28 multi_7x28_mod_11907(clk,rst,matrix_A[11907],matrix_B[107],mul_res1[11907]);
multi_7x28 multi_7x28_mod_11908(clk,rst,matrix_A[11908],matrix_B[108],mul_res1[11908]);
multi_7x28 multi_7x28_mod_11909(clk,rst,matrix_A[11909],matrix_B[109],mul_res1[11909]);
multi_7x28 multi_7x28_mod_11910(clk,rst,matrix_A[11910],matrix_B[110],mul_res1[11910]);
multi_7x28 multi_7x28_mod_11911(clk,rst,matrix_A[11911],matrix_B[111],mul_res1[11911]);
multi_7x28 multi_7x28_mod_11912(clk,rst,matrix_A[11912],matrix_B[112],mul_res1[11912]);
multi_7x28 multi_7x28_mod_11913(clk,rst,matrix_A[11913],matrix_B[113],mul_res1[11913]);
multi_7x28 multi_7x28_mod_11914(clk,rst,matrix_A[11914],matrix_B[114],mul_res1[11914]);
multi_7x28 multi_7x28_mod_11915(clk,rst,matrix_A[11915],matrix_B[115],mul_res1[11915]);
multi_7x28 multi_7x28_mod_11916(clk,rst,matrix_A[11916],matrix_B[116],mul_res1[11916]);
multi_7x28 multi_7x28_mod_11917(clk,rst,matrix_A[11917],matrix_B[117],mul_res1[11917]);
multi_7x28 multi_7x28_mod_11918(clk,rst,matrix_A[11918],matrix_B[118],mul_res1[11918]);
multi_7x28 multi_7x28_mod_11919(clk,rst,matrix_A[11919],matrix_B[119],mul_res1[11919]);
multi_7x28 multi_7x28_mod_11920(clk,rst,matrix_A[11920],matrix_B[120],mul_res1[11920]);
multi_7x28 multi_7x28_mod_11921(clk,rst,matrix_A[11921],matrix_B[121],mul_res1[11921]);
multi_7x28 multi_7x28_mod_11922(clk,rst,matrix_A[11922],matrix_B[122],mul_res1[11922]);
multi_7x28 multi_7x28_mod_11923(clk,rst,matrix_A[11923],matrix_B[123],mul_res1[11923]);
multi_7x28 multi_7x28_mod_11924(clk,rst,matrix_A[11924],matrix_B[124],mul_res1[11924]);
multi_7x28 multi_7x28_mod_11925(clk,rst,matrix_A[11925],matrix_B[125],mul_res1[11925]);
multi_7x28 multi_7x28_mod_11926(clk,rst,matrix_A[11926],matrix_B[126],mul_res1[11926]);
multi_7x28 multi_7x28_mod_11927(clk,rst,matrix_A[11927],matrix_B[127],mul_res1[11927]);
multi_7x28 multi_7x28_mod_11928(clk,rst,matrix_A[11928],matrix_B[128],mul_res1[11928]);
multi_7x28 multi_7x28_mod_11929(clk,rst,matrix_A[11929],matrix_B[129],mul_res1[11929]);
multi_7x28 multi_7x28_mod_11930(clk,rst,matrix_A[11930],matrix_B[130],mul_res1[11930]);
multi_7x28 multi_7x28_mod_11931(clk,rst,matrix_A[11931],matrix_B[131],mul_res1[11931]);
multi_7x28 multi_7x28_mod_11932(clk,rst,matrix_A[11932],matrix_B[132],mul_res1[11932]);
multi_7x28 multi_7x28_mod_11933(clk,rst,matrix_A[11933],matrix_B[133],mul_res1[11933]);
multi_7x28 multi_7x28_mod_11934(clk,rst,matrix_A[11934],matrix_B[134],mul_res1[11934]);
multi_7x28 multi_7x28_mod_11935(clk,rst,matrix_A[11935],matrix_B[135],mul_res1[11935]);
multi_7x28 multi_7x28_mod_11936(clk,rst,matrix_A[11936],matrix_B[136],mul_res1[11936]);
multi_7x28 multi_7x28_mod_11937(clk,rst,matrix_A[11937],matrix_B[137],mul_res1[11937]);
multi_7x28 multi_7x28_mod_11938(clk,rst,matrix_A[11938],matrix_B[138],mul_res1[11938]);
multi_7x28 multi_7x28_mod_11939(clk,rst,matrix_A[11939],matrix_B[139],mul_res1[11939]);
multi_7x28 multi_7x28_mod_11940(clk,rst,matrix_A[11940],matrix_B[140],mul_res1[11940]);
multi_7x28 multi_7x28_mod_11941(clk,rst,matrix_A[11941],matrix_B[141],mul_res1[11941]);
multi_7x28 multi_7x28_mod_11942(clk,rst,matrix_A[11942],matrix_B[142],mul_res1[11942]);
multi_7x28 multi_7x28_mod_11943(clk,rst,matrix_A[11943],matrix_B[143],mul_res1[11943]);
multi_7x28 multi_7x28_mod_11944(clk,rst,matrix_A[11944],matrix_B[144],mul_res1[11944]);
multi_7x28 multi_7x28_mod_11945(clk,rst,matrix_A[11945],matrix_B[145],mul_res1[11945]);
multi_7x28 multi_7x28_mod_11946(clk,rst,matrix_A[11946],matrix_B[146],mul_res1[11946]);
multi_7x28 multi_7x28_mod_11947(clk,rst,matrix_A[11947],matrix_B[147],mul_res1[11947]);
multi_7x28 multi_7x28_mod_11948(clk,rst,matrix_A[11948],matrix_B[148],mul_res1[11948]);
multi_7x28 multi_7x28_mod_11949(clk,rst,matrix_A[11949],matrix_B[149],mul_res1[11949]);
multi_7x28 multi_7x28_mod_11950(clk,rst,matrix_A[11950],matrix_B[150],mul_res1[11950]);
multi_7x28 multi_7x28_mod_11951(clk,rst,matrix_A[11951],matrix_B[151],mul_res1[11951]);
multi_7x28 multi_7x28_mod_11952(clk,rst,matrix_A[11952],matrix_B[152],mul_res1[11952]);
multi_7x28 multi_7x28_mod_11953(clk,rst,matrix_A[11953],matrix_B[153],mul_res1[11953]);
multi_7x28 multi_7x28_mod_11954(clk,rst,matrix_A[11954],matrix_B[154],mul_res1[11954]);
multi_7x28 multi_7x28_mod_11955(clk,rst,matrix_A[11955],matrix_B[155],mul_res1[11955]);
multi_7x28 multi_7x28_mod_11956(clk,rst,matrix_A[11956],matrix_B[156],mul_res1[11956]);
multi_7x28 multi_7x28_mod_11957(clk,rst,matrix_A[11957],matrix_B[157],mul_res1[11957]);
multi_7x28 multi_7x28_mod_11958(clk,rst,matrix_A[11958],matrix_B[158],mul_res1[11958]);
multi_7x28 multi_7x28_mod_11959(clk,rst,matrix_A[11959],matrix_B[159],mul_res1[11959]);
multi_7x28 multi_7x28_mod_11960(clk,rst,matrix_A[11960],matrix_B[160],mul_res1[11960]);
multi_7x28 multi_7x28_mod_11961(clk,rst,matrix_A[11961],matrix_B[161],mul_res1[11961]);
multi_7x28 multi_7x28_mod_11962(clk,rst,matrix_A[11962],matrix_B[162],mul_res1[11962]);
multi_7x28 multi_7x28_mod_11963(clk,rst,matrix_A[11963],matrix_B[163],mul_res1[11963]);
multi_7x28 multi_7x28_mod_11964(clk,rst,matrix_A[11964],matrix_B[164],mul_res1[11964]);
multi_7x28 multi_7x28_mod_11965(clk,rst,matrix_A[11965],matrix_B[165],mul_res1[11965]);
multi_7x28 multi_7x28_mod_11966(clk,rst,matrix_A[11966],matrix_B[166],mul_res1[11966]);
multi_7x28 multi_7x28_mod_11967(clk,rst,matrix_A[11967],matrix_B[167],mul_res1[11967]);
multi_7x28 multi_7x28_mod_11968(clk,rst,matrix_A[11968],matrix_B[168],mul_res1[11968]);
multi_7x28 multi_7x28_mod_11969(clk,rst,matrix_A[11969],matrix_B[169],mul_res1[11969]);
multi_7x28 multi_7x28_mod_11970(clk,rst,matrix_A[11970],matrix_B[170],mul_res1[11970]);
multi_7x28 multi_7x28_mod_11971(clk,rst,matrix_A[11971],matrix_B[171],mul_res1[11971]);
multi_7x28 multi_7x28_mod_11972(clk,rst,matrix_A[11972],matrix_B[172],mul_res1[11972]);
multi_7x28 multi_7x28_mod_11973(clk,rst,matrix_A[11973],matrix_B[173],mul_res1[11973]);
multi_7x28 multi_7x28_mod_11974(clk,rst,matrix_A[11974],matrix_B[174],mul_res1[11974]);
multi_7x28 multi_7x28_mod_11975(clk,rst,matrix_A[11975],matrix_B[175],mul_res1[11975]);
multi_7x28 multi_7x28_mod_11976(clk,rst,matrix_A[11976],matrix_B[176],mul_res1[11976]);
multi_7x28 multi_7x28_mod_11977(clk,rst,matrix_A[11977],matrix_B[177],mul_res1[11977]);
multi_7x28 multi_7x28_mod_11978(clk,rst,matrix_A[11978],matrix_B[178],mul_res1[11978]);
multi_7x28 multi_7x28_mod_11979(clk,rst,matrix_A[11979],matrix_B[179],mul_res1[11979]);
multi_7x28 multi_7x28_mod_11980(clk,rst,matrix_A[11980],matrix_B[180],mul_res1[11980]);
multi_7x28 multi_7x28_mod_11981(clk,rst,matrix_A[11981],matrix_B[181],mul_res1[11981]);
multi_7x28 multi_7x28_mod_11982(clk,rst,matrix_A[11982],matrix_B[182],mul_res1[11982]);
multi_7x28 multi_7x28_mod_11983(clk,rst,matrix_A[11983],matrix_B[183],mul_res1[11983]);
multi_7x28 multi_7x28_mod_11984(clk,rst,matrix_A[11984],matrix_B[184],mul_res1[11984]);
multi_7x28 multi_7x28_mod_11985(clk,rst,matrix_A[11985],matrix_B[185],mul_res1[11985]);
multi_7x28 multi_7x28_mod_11986(clk,rst,matrix_A[11986],matrix_B[186],mul_res1[11986]);
multi_7x28 multi_7x28_mod_11987(clk,rst,matrix_A[11987],matrix_B[187],mul_res1[11987]);
multi_7x28 multi_7x28_mod_11988(clk,rst,matrix_A[11988],matrix_B[188],mul_res1[11988]);
multi_7x28 multi_7x28_mod_11989(clk,rst,matrix_A[11989],matrix_B[189],mul_res1[11989]);
multi_7x28 multi_7x28_mod_11990(clk,rst,matrix_A[11990],matrix_B[190],mul_res1[11990]);
multi_7x28 multi_7x28_mod_11991(clk,rst,matrix_A[11991],matrix_B[191],mul_res1[11991]);
multi_7x28 multi_7x28_mod_11992(clk,rst,matrix_A[11992],matrix_B[192],mul_res1[11992]);
multi_7x28 multi_7x28_mod_11993(clk,rst,matrix_A[11993],matrix_B[193],mul_res1[11993]);
multi_7x28 multi_7x28_mod_11994(clk,rst,matrix_A[11994],matrix_B[194],mul_res1[11994]);
multi_7x28 multi_7x28_mod_11995(clk,rst,matrix_A[11995],matrix_B[195],mul_res1[11995]);
multi_7x28 multi_7x28_mod_11996(clk,rst,matrix_A[11996],matrix_B[196],mul_res1[11996]);
multi_7x28 multi_7x28_mod_11997(clk,rst,matrix_A[11997],matrix_B[197],mul_res1[11997]);
multi_7x28 multi_7x28_mod_11998(clk,rst,matrix_A[11998],matrix_B[198],mul_res1[11998]);
multi_7x28 multi_7x28_mod_11999(clk,rst,matrix_A[11999],matrix_B[199],mul_res1[11999]);
multi_7x28 multi_7x28_mod_12000(clk,rst,matrix_A[12000],matrix_B[0],mul_res1[12000]);
multi_7x28 multi_7x28_mod_12001(clk,rst,matrix_A[12001],matrix_B[1],mul_res1[12001]);
multi_7x28 multi_7x28_mod_12002(clk,rst,matrix_A[12002],matrix_B[2],mul_res1[12002]);
multi_7x28 multi_7x28_mod_12003(clk,rst,matrix_A[12003],matrix_B[3],mul_res1[12003]);
multi_7x28 multi_7x28_mod_12004(clk,rst,matrix_A[12004],matrix_B[4],mul_res1[12004]);
multi_7x28 multi_7x28_mod_12005(clk,rst,matrix_A[12005],matrix_B[5],mul_res1[12005]);
multi_7x28 multi_7x28_mod_12006(clk,rst,matrix_A[12006],matrix_B[6],mul_res1[12006]);
multi_7x28 multi_7x28_mod_12007(clk,rst,matrix_A[12007],matrix_B[7],mul_res1[12007]);
multi_7x28 multi_7x28_mod_12008(clk,rst,matrix_A[12008],matrix_B[8],mul_res1[12008]);
multi_7x28 multi_7x28_mod_12009(clk,rst,matrix_A[12009],matrix_B[9],mul_res1[12009]);
multi_7x28 multi_7x28_mod_12010(clk,rst,matrix_A[12010],matrix_B[10],mul_res1[12010]);
multi_7x28 multi_7x28_mod_12011(clk,rst,matrix_A[12011],matrix_B[11],mul_res1[12011]);
multi_7x28 multi_7x28_mod_12012(clk,rst,matrix_A[12012],matrix_B[12],mul_res1[12012]);
multi_7x28 multi_7x28_mod_12013(clk,rst,matrix_A[12013],matrix_B[13],mul_res1[12013]);
multi_7x28 multi_7x28_mod_12014(clk,rst,matrix_A[12014],matrix_B[14],mul_res1[12014]);
multi_7x28 multi_7x28_mod_12015(clk,rst,matrix_A[12015],matrix_B[15],mul_res1[12015]);
multi_7x28 multi_7x28_mod_12016(clk,rst,matrix_A[12016],matrix_B[16],mul_res1[12016]);
multi_7x28 multi_7x28_mod_12017(clk,rst,matrix_A[12017],matrix_B[17],mul_res1[12017]);
multi_7x28 multi_7x28_mod_12018(clk,rst,matrix_A[12018],matrix_B[18],mul_res1[12018]);
multi_7x28 multi_7x28_mod_12019(clk,rst,matrix_A[12019],matrix_B[19],mul_res1[12019]);
multi_7x28 multi_7x28_mod_12020(clk,rst,matrix_A[12020],matrix_B[20],mul_res1[12020]);
multi_7x28 multi_7x28_mod_12021(clk,rst,matrix_A[12021],matrix_B[21],mul_res1[12021]);
multi_7x28 multi_7x28_mod_12022(clk,rst,matrix_A[12022],matrix_B[22],mul_res1[12022]);
multi_7x28 multi_7x28_mod_12023(clk,rst,matrix_A[12023],matrix_B[23],mul_res1[12023]);
multi_7x28 multi_7x28_mod_12024(clk,rst,matrix_A[12024],matrix_B[24],mul_res1[12024]);
multi_7x28 multi_7x28_mod_12025(clk,rst,matrix_A[12025],matrix_B[25],mul_res1[12025]);
multi_7x28 multi_7x28_mod_12026(clk,rst,matrix_A[12026],matrix_B[26],mul_res1[12026]);
multi_7x28 multi_7x28_mod_12027(clk,rst,matrix_A[12027],matrix_B[27],mul_res1[12027]);
multi_7x28 multi_7x28_mod_12028(clk,rst,matrix_A[12028],matrix_B[28],mul_res1[12028]);
multi_7x28 multi_7x28_mod_12029(clk,rst,matrix_A[12029],matrix_B[29],mul_res1[12029]);
multi_7x28 multi_7x28_mod_12030(clk,rst,matrix_A[12030],matrix_B[30],mul_res1[12030]);
multi_7x28 multi_7x28_mod_12031(clk,rst,matrix_A[12031],matrix_B[31],mul_res1[12031]);
multi_7x28 multi_7x28_mod_12032(clk,rst,matrix_A[12032],matrix_B[32],mul_res1[12032]);
multi_7x28 multi_7x28_mod_12033(clk,rst,matrix_A[12033],matrix_B[33],mul_res1[12033]);
multi_7x28 multi_7x28_mod_12034(clk,rst,matrix_A[12034],matrix_B[34],mul_res1[12034]);
multi_7x28 multi_7x28_mod_12035(clk,rst,matrix_A[12035],matrix_B[35],mul_res1[12035]);
multi_7x28 multi_7x28_mod_12036(clk,rst,matrix_A[12036],matrix_B[36],mul_res1[12036]);
multi_7x28 multi_7x28_mod_12037(clk,rst,matrix_A[12037],matrix_B[37],mul_res1[12037]);
multi_7x28 multi_7x28_mod_12038(clk,rst,matrix_A[12038],matrix_B[38],mul_res1[12038]);
multi_7x28 multi_7x28_mod_12039(clk,rst,matrix_A[12039],matrix_B[39],mul_res1[12039]);
multi_7x28 multi_7x28_mod_12040(clk,rst,matrix_A[12040],matrix_B[40],mul_res1[12040]);
multi_7x28 multi_7x28_mod_12041(clk,rst,matrix_A[12041],matrix_B[41],mul_res1[12041]);
multi_7x28 multi_7x28_mod_12042(clk,rst,matrix_A[12042],matrix_B[42],mul_res1[12042]);
multi_7x28 multi_7x28_mod_12043(clk,rst,matrix_A[12043],matrix_B[43],mul_res1[12043]);
multi_7x28 multi_7x28_mod_12044(clk,rst,matrix_A[12044],matrix_B[44],mul_res1[12044]);
multi_7x28 multi_7x28_mod_12045(clk,rst,matrix_A[12045],matrix_B[45],mul_res1[12045]);
multi_7x28 multi_7x28_mod_12046(clk,rst,matrix_A[12046],matrix_B[46],mul_res1[12046]);
multi_7x28 multi_7x28_mod_12047(clk,rst,matrix_A[12047],matrix_B[47],mul_res1[12047]);
multi_7x28 multi_7x28_mod_12048(clk,rst,matrix_A[12048],matrix_B[48],mul_res1[12048]);
multi_7x28 multi_7x28_mod_12049(clk,rst,matrix_A[12049],matrix_B[49],mul_res1[12049]);
multi_7x28 multi_7x28_mod_12050(clk,rst,matrix_A[12050],matrix_B[50],mul_res1[12050]);
multi_7x28 multi_7x28_mod_12051(clk,rst,matrix_A[12051],matrix_B[51],mul_res1[12051]);
multi_7x28 multi_7x28_mod_12052(clk,rst,matrix_A[12052],matrix_B[52],mul_res1[12052]);
multi_7x28 multi_7x28_mod_12053(clk,rst,matrix_A[12053],matrix_B[53],mul_res1[12053]);
multi_7x28 multi_7x28_mod_12054(clk,rst,matrix_A[12054],matrix_B[54],mul_res1[12054]);
multi_7x28 multi_7x28_mod_12055(clk,rst,matrix_A[12055],matrix_B[55],mul_res1[12055]);
multi_7x28 multi_7x28_mod_12056(clk,rst,matrix_A[12056],matrix_B[56],mul_res1[12056]);
multi_7x28 multi_7x28_mod_12057(clk,rst,matrix_A[12057],matrix_B[57],mul_res1[12057]);
multi_7x28 multi_7x28_mod_12058(clk,rst,matrix_A[12058],matrix_B[58],mul_res1[12058]);
multi_7x28 multi_7x28_mod_12059(clk,rst,matrix_A[12059],matrix_B[59],mul_res1[12059]);
multi_7x28 multi_7x28_mod_12060(clk,rst,matrix_A[12060],matrix_B[60],mul_res1[12060]);
multi_7x28 multi_7x28_mod_12061(clk,rst,matrix_A[12061],matrix_B[61],mul_res1[12061]);
multi_7x28 multi_7x28_mod_12062(clk,rst,matrix_A[12062],matrix_B[62],mul_res1[12062]);
multi_7x28 multi_7x28_mod_12063(clk,rst,matrix_A[12063],matrix_B[63],mul_res1[12063]);
multi_7x28 multi_7x28_mod_12064(clk,rst,matrix_A[12064],matrix_B[64],mul_res1[12064]);
multi_7x28 multi_7x28_mod_12065(clk,rst,matrix_A[12065],matrix_B[65],mul_res1[12065]);
multi_7x28 multi_7x28_mod_12066(clk,rst,matrix_A[12066],matrix_B[66],mul_res1[12066]);
multi_7x28 multi_7x28_mod_12067(clk,rst,matrix_A[12067],matrix_B[67],mul_res1[12067]);
multi_7x28 multi_7x28_mod_12068(clk,rst,matrix_A[12068],matrix_B[68],mul_res1[12068]);
multi_7x28 multi_7x28_mod_12069(clk,rst,matrix_A[12069],matrix_B[69],mul_res1[12069]);
multi_7x28 multi_7x28_mod_12070(clk,rst,matrix_A[12070],matrix_B[70],mul_res1[12070]);
multi_7x28 multi_7x28_mod_12071(clk,rst,matrix_A[12071],matrix_B[71],mul_res1[12071]);
multi_7x28 multi_7x28_mod_12072(clk,rst,matrix_A[12072],matrix_B[72],mul_res1[12072]);
multi_7x28 multi_7x28_mod_12073(clk,rst,matrix_A[12073],matrix_B[73],mul_res1[12073]);
multi_7x28 multi_7x28_mod_12074(clk,rst,matrix_A[12074],matrix_B[74],mul_res1[12074]);
multi_7x28 multi_7x28_mod_12075(clk,rst,matrix_A[12075],matrix_B[75],mul_res1[12075]);
multi_7x28 multi_7x28_mod_12076(clk,rst,matrix_A[12076],matrix_B[76],mul_res1[12076]);
multi_7x28 multi_7x28_mod_12077(clk,rst,matrix_A[12077],matrix_B[77],mul_res1[12077]);
multi_7x28 multi_7x28_mod_12078(clk,rst,matrix_A[12078],matrix_B[78],mul_res1[12078]);
multi_7x28 multi_7x28_mod_12079(clk,rst,matrix_A[12079],matrix_B[79],mul_res1[12079]);
multi_7x28 multi_7x28_mod_12080(clk,rst,matrix_A[12080],matrix_B[80],mul_res1[12080]);
multi_7x28 multi_7x28_mod_12081(clk,rst,matrix_A[12081],matrix_B[81],mul_res1[12081]);
multi_7x28 multi_7x28_mod_12082(clk,rst,matrix_A[12082],matrix_B[82],mul_res1[12082]);
multi_7x28 multi_7x28_mod_12083(clk,rst,matrix_A[12083],matrix_B[83],mul_res1[12083]);
multi_7x28 multi_7x28_mod_12084(clk,rst,matrix_A[12084],matrix_B[84],mul_res1[12084]);
multi_7x28 multi_7x28_mod_12085(clk,rst,matrix_A[12085],matrix_B[85],mul_res1[12085]);
multi_7x28 multi_7x28_mod_12086(clk,rst,matrix_A[12086],matrix_B[86],mul_res1[12086]);
multi_7x28 multi_7x28_mod_12087(clk,rst,matrix_A[12087],matrix_B[87],mul_res1[12087]);
multi_7x28 multi_7x28_mod_12088(clk,rst,matrix_A[12088],matrix_B[88],mul_res1[12088]);
multi_7x28 multi_7x28_mod_12089(clk,rst,matrix_A[12089],matrix_B[89],mul_res1[12089]);
multi_7x28 multi_7x28_mod_12090(clk,rst,matrix_A[12090],matrix_B[90],mul_res1[12090]);
multi_7x28 multi_7x28_mod_12091(clk,rst,matrix_A[12091],matrix_B[91],mul_res1[12091]);
multi_7x28 multi_7x28_mod_12092(clk,rst,matrix_A[12092],matrix_B[92],mul_res1[12092]);
multi_7x28 multi_7x28_mod_12093(clk,rst,matrix_A[12093],matrix_B[93],mul_res1[12093]);
multi_7x28 multi_7x28_mod_12094(clk,rst,matrix_A[12094],matrix_B[94],mul_res1[12094]);
multi_7x28 multi_7x28_mod_12095(clk,rst,matrix_A[12095],matrix_B[95],mul_res1[12095]);
multi_7x28 multi_7x28_mod_12096(clk,rst,matrix_A[12096],matrix_B[96],mul_res1[12096]);
multi_7x28 multi_7x28_mod_12097(clk,rst,matrix_A[12097],matrix_B[97],mul_res1[12097]);
multi_7x28 multi_7x28_mod_12098(clk,rst,matrix_A[12098],matrix_B[98],mul_res1[12098]);
multi_7x28 multi_7x28_mod_12099(clk,rst,matrix_A[12099],matrix_B[99],mul_res1[12099]);
multi_7x28 multi_7x28_mod_12100(clk,rst,matrix_A[12100],matrix_B[100],mul_res1[12100]);
multi_7x28 multi_7x28_mod_12101(clk,rst,matrix_A[12101],matrix_B[101],mul_res1[12101]);
multi_7x28 multi_7x28_mod_12102(clk,rst,matrix_A[12102],matrix_B[102],mul_res1[12102]);
multi_7x28 multi_7x28_mod_12103(clk,rst,matrix_A[12103],matrix_B[103],mul_res1[12103]);
multi_7x28 multi_7x28_mod_12104(clk,rst,matrix_A[12104],matrix_B[104],mul_res1[12104]);
multi_7x28 multi_7x28_mod_12105(clk,rst,matrix_A[12105],matrix_B[105],mul_res1[12105]);
multi_7x28 multi_7x28_mod_12106(clk,rst,matrix_A[12106],matrix_B[106],mul_res1[12106]);
multi_7x28 multi_7x28_mod_12107(clk,rst,matrix_A[12107],matrix_B[107],mul_res1[12107]);
multi_7x28 multi_7x28_mod_12108(clk,rst,matrix_A[12108],matrix_B[108],mul_res1[12108]);
multi_7x28 multi_7x28_mod_12109(clk,rst,matrix_A[12109],matrix_B[109],mul_res1[12109]);
multi_7x28 multi_7x28_mod_12110(clk,rst,matrix_A[12110],matrix_B[110],mul_res1[12110]);
multi_7x28 multi_7x28_mod_12111(clk,rst,matrix_A[12111],matrix_B[111],mul_res1[12111]);
multi_7x28 multi_7x28_mod_12112(clk,rst,matrix_A[12112],matrix_B[112],mul_res1[12112]);
multi_7x28 multi_7x28_mod_12113(clk,rst,matrix_A[12113],matrix_B[113],mul_res1[12113]);
multi_7x28 multi_7x28_mod_12114(clk,rst,matrix_A[12114],matrix_B[114],mul_res1[12114]);
multi_7x28 multi_7x28_mod_12115(clk,rst,matrix_A[12115],matrix_B[115],mul_res1[12115]);
multi_7x28 multi_7x28_mod_12116(clk,rst,matrix_A[12116],matrix_B[116],mul_res1[12116]);
multi_7x28 multi_7x28_mod_12117(clk,rst,matrix_A[12117],matrix_B[117],mul_res1[12117]);
multi_7x28 multi_7x28_mod_12118(clk,rst,matrix_A[12118],matrix_B[118],mul_res1[12118]);
multi_7x28 multi_7x28_mod_12119(clk,rst,matrix_A[12119],matrix_B[119],mul_res1[12119]);
multi_7x28 multi_7x28_mod_12120(clk,rst,matrix_A[12120],matrix_B[120],mul_res1[12120]);
multi_7x28 multi_7x28_mod_12121(clk,rst,matrix_A[12121],matrix_B[121],mul_res1[12121]);
multi_7x28 multi_7x28_mod_12122(clk,rst,matrix_A[12122],matrix_B[122],mul_res1[12122]);
multi_7x28 multi_7x28_mod_12123(clk,rst,matrix_A[12123],matrix_B[123],mul_res1[12123]);
multi_7x28 multi_7x28_mod_12124(clk,rst,matrix_A[12124],matrix_B[124],mul_res1[12124]);
multi_7x28 multi_7x28_mod_12125(clk,rst,matrix_A[12125],matrix_B[125],mul_res1[12125]);
multi_7x28 multi_7x28_mod_12126(clk,rst,matrix_A[12126],matrix_B[126],mul_res1[12126]);
multi_7x28 multi_7x28_mod_12127(clk,rst,matrix_A[12127],matrix_B[127],mul_res1[12127]);
multi_7x28 multi_7x28_mod_12128(clk,rst,matrix_A[12128],matrix_B[128],mul_res1[12128]);
multi_7x28 multi_7x28_mod_12129(clk,rst,matrix_A[12129],matrix_B[129],mul_res1[12129]);
multi_7x28 multi_7x28_mod_12130(clk,rst,matrix_A[12130],matrix_B[130],mul_res1[12130]);
multi_7x28 multi_7x28_mod_12131(clk,rst,matrix_A[12131],matrix_B[131],mul_res1[12131]);
multi_7x28 multi_7x28_mod_12132(clk,rst,matrix_A[12132],matrix_B[132],mul_res1[12132]);
multi_7x28 multi_7x28_mod_12133(clk,rst,matrix_A[12133],matrix_B[133],mul_res1[12133]);
multi_7x28 multi_7x28_mod_12134(clk,rst,matrix_A[12134],matrix_B[134],mul_res1[12134]);
multi_7x28 multi_7x28_mod_12135(clk,rst,matrix_A[12135],matrix_B[135],mul_res1[12135]);
multi_7x28 multi_7x28_mod_12136(clk,rst,matrix_A[12136],matrix_B[136],mul_res1[12136]);
multi_7x28 multi_7x28_mod_12137(clk,rst,matrix_A[12137],matrix_B[137],mul_res1[12137]);
multi_7x28 multi_7x28_mod_12138(clk,rst,matrix_A[12138],matrix_B[138],mul_res1[12138]);
multi_7x28 multi_7x28_mod_12139(clk,rst,matrix_A[12139],matrix_B[139],mul_res1[12139]);
multi_7x28 multi_7x28_mod_12140(clk,rst,matrix_A[12140],matrix_B[140],mul_res1[12140]);
multi_7x28 multi_7x28_mod_12141(clk,rst,matrix_A[12141],matrix_B[141],mul_res1[12141]);
multi_7x28 multi_7x28_mod_12142(clk,rst,matrix_A[12142],matrix_B[142],mul_res1[12142]);
multi_7x28 multi_7x28_mod_12143(clk,rst,matrix_A[12143],matrix_B[143],mul_res1[12143]);
multi_7x28 multi_7x28_mod_12144(clk,rst,matrix_A[12144],matrix_B[144],mul_res1[12144]);
multi_7x28 multi_7x28_mod_12145(clk,rst,matrix_A[12145],matrix_B[145],mul_res1[12145]);
multi_7x28 multi_7x28_mod_12146(clk,rst,matrix_A[12146],matrix_B[146],mul_res1[12146]);
multi_7x28 multi_7x28_mod_12147(clk,rst,matrix_A[12147],matrix_B[147],mul_res1[12147]);
multi_7x28 multi_7x28_mod_12148(clk,rst,matrix_A[12148],matrix_B[148],mul_res1[12148]);
multi_7x28 multi_7x28_mod_12149(clk,rst,matrix_A[12149],matrix_B[149],mul_res1[12149]);
multi_7x28 multi_7x28_mod_12150(clk,rst,matrix_A[12150],matrix_B[150],mul_res1[12150]);
multi_7x28 multi_7x28_mod_12151(clk,rst,matrix_A[12151],matrix_B[151],mul_res1[12151]);
multi_7x28 multi_7x28_mod_12152(clk,rst,matrix_A[12152],matrix_B[152],mul_res1[12152]);
multi_7x28 multi_7x28_mod_12153(clk,rst,matrix_A[12153],matrix_B[153],mul_res1[12153]);
multi_7x28 multi_7x28_mod_12154(clk,rst,matrix_A[12154],matrix_B[154],mul_res1[12154]);
multi_7x28 multi_7x28_mod_12155(clk,rst,matrix_A[12155],matrix_B[155],mul_res1[12155]);
multi_7x28 multi_7x28_mod_12156(clk,rst,matrix_A[12156],matrix_B[156],mul_res1[12156]);
multi_7x28 multi_7x28_mod_12157(clk,rst,matrix_A[12157],matrix_B[157],mul_res1[12157]);
multi_7x28 multi_7x28_mod_12158(clk,rst,matrix_A[12158],matrix_B[158],mul_res1[12158]);
multi_7x28 multi_7x28_mod_12159(clk,rst,matrix_A[12159],matrix_B[159],mul_res1[12159]);
multi_7x28 multi_7x28_mod_12160(clk,rst,matrix_A[12160],matrix_B[160],mul_res1[12160]);
multi_7x28 multi_7x28_mod_12161(clk,rst,matrix_A[12161],matrix_B[161],mul_res1[12161]);
multi_7x28 multi_7x28_mod_12162(clk,rst,matrix_A[12162],matrix_B[162],mul_res1[12162]);
multi_7x28 multi_7x28_mod_12163(clk,rst,matrix_A[12163],matrix_B[163],mul_res1[12163]);
multi_7x28 multi_7x28_mod_12164(clk,rst,matrix_A[12164],matrix_B[164],mul_res1[12164]);
multi_7x28 multi_7x28_mod_12165(clk,rst,matrix_A[12165],matrix_B[165],mul_res1[12165]);
multi_7x28 multi_7x28_mod_12166(clk,rst,matrix_A[12166],matrix_B[166],mul_res1[12166]);
multi_7x28 multi_7x28_mod_12167(clk,rst,matrix_A[12167],matrix_B[167],mul_res1[12167]);
multi_7x28 multi_7x28_mod_12168(clk,rst,matrix_A[12168],matrix_B[168],mul_res1[12168]);
multi_7x28 multi_7x28_mod_12169(clk,rst,matrix_A[12169],matrix_B[169],mul_res1[12169]);
multi_7x28 multi_7x28_mod_12170(clk,rst,matrix_A[12170],matrix_B[170],mul_res1[12170]);
multi_7x28 multi_7x28_mod_12171(clk,rst,matrix_A[12171],matrix_B[171],mul_res1[12171]);
multi_7x28 multi_7x28_mod_12172(clk,rst,matrix_A[12172],matrix_B[172],mul_res1[12172]);
multi_7x28 multi_7x28_mod_12173(clk,rst,matrix_A[12173],matrix_B[173],mul_res1[12173]);
multi_7x28 multi_7x28_mod_12174(clk,rst,matrix_A[12174],matrix_B[174],mul_res1[12174]);
multi_7x28 multi_7x28_mod_12175(clk,rst,matrix_A[12175],matrix_B[175],mul_res1[12175]);
multi_7x28 multi_7x28_mod_12176(clk,rst,matrix_A[12176],matrix_B[176],mul_res1[12176]);
multi_7x28 multi_7x28_mod_12177(clk,rst,matrix_A[12177],matrix_B[177],mul_res1[12177]);
multi_7x28 multi_7x28_mod_12178(clk,rst,matrix_A[12178],matrix_B[178],mul_res1[12178]);
multi_7x28 multi_7x28_mod_12179(clk,rst,matrix_A[12179],matrix_B[179],mul_res1[12179]);
multi_7x28 multi_7x28_mod_12180(clk,rst,matrix_A[12180],matrix_B[180],mul_res1[12180]);
multi_7x28 multi_7x28_mod_12181(clk,rst,matrix_A[12181],matrix_B[181],mul_res1[12181]);
multi_7x28 multi_7x28_mod_12182(clk,rst,matrix_A[12182],matrix_B[182],mul_res1[12182]);
multi_7x28 multi_7x28_mod_12183(clk,rst,matrix_A[12183],matrix_B[183],mul_res1[12183]);
multi_7x28 multi_7x28_mod_12184(clk,rst,matrix_A[12184],matrix_B[184],mul_res1[12184]);
multi_7x28 multi_7x28_mod_12185(clk,rst,matrix_A[12185],matrix_B[185],mul_res1[12185]);
multi_7x28 multi_7x28_mod_12186(clk,rst,matrix_A[12186],matrix_B[186],mul_res1[12186]);
multi_7x28 multi_7x28_mod_12187(clk,rst,matrix_A[12187],matrix_B[187],mul_res1[12187]);
multi_7x28 multi_7x28_mod_12188(clk,rst,matrix_A[12188],matrix_B[188],mul_res1[12188]);
multi_7x28 multi_7x28_mod_12189(clk,rst,matrix_A[12189],matrix_B[189],mul_res1[12189]);
multi_7x28 multi_7x28_mod_12190(clk,rst,matrix_A[12190],matrix_B[190],mul_res1[12190]);
multi_7x28 multi_7x28_mod_12191(clk,rst,matrix_A[12191],matrix_B[191],mul_res1[12191]);
multi_7x28 multi_7x28_mod_12192(clk,rst,matrix_A[12192],matrix_B[192],mul_res1[12192]);
multi_7x28 multi_7x28_mod_12193(clk,rst,matrix_A[12193],matrix_B[193],mul_res1[12193]);
multi_7x28 multi_7x28_mod_12194(clk,rst,matrix_A[12194],matrix_B[194],mul_res1[12194]);
multi_7x28 multi_7x28_mod_12195(clk,rst,matrix_A[12195],matrix_B[195],mul_res1[12195]);
multi_7x28 multi_7x28_mod_12196(clk,rst,matrix_A[12196],matrix_B[196],mul_res1[12196]);
multi_7x28 multi_7x28_mod_12197(clk,rst,matrix_A[12197],matrix_B[197],mul_res1[12197]);
multi_7x28 multi_7x28_mod_12198(clk,rst,matrix_A[12198],matrix_B[198],mul_res1[12198]);
multi_7x28 multi_7x28_mod_12199(clk,rst,matrix_A[12199],matrix_B[199],mul_res1[12199]);
multi_7x28 multi_7x28_mod_12200(clk,rst,matrix_A[12200],matrix_B[0],mul_res1[12200]);
multi_7x28 multi_7x28_mod_12201(clk,rst,matrix_A[12201],matrix_B[1],mul_res1[12201]);
multi_7x28 multi_7x28_mod_12202(clk,rst,matrix_A[12202],matrix_B[2],mul_res1[12202]);
multi_7x28 multi_7x28_mod_12203(clk,rst,matrix_A[12203],matrix_B[3],mul_res1[12203]);
multi_7x28 multi_7x28_mod_12204(clk,rst,matrix_A[12204],matrix_B[4],mul_res1[12204]);
multi_7x28 multi_7x28_mod_12205(clk,rst,matrix_A[12205],matrix_B[5],mul_res1[12205]);
multi_7x28 multi_7x28_mod_12206(clk,rst,matrix_A[12206],matrix_B[6],mul_res1[12206]);
multi_7x28 multi_7x28_mod_12207(clk,rst,matrix_A[12207],matrix_B[7],mul_res1[12207]);
multi_7x28 multi_7x28_mod_12208(clk,rst,matrix_A[12208],matrix_B[8],mul_res1[12208]);
multi_7x28 multi_7x28_mod_12209(clk,rst,matrix_A[12209],matrix_B[9],mul_res1[12209]);
multi_7x28 multi_7x28_mod_12210(clk,rst,matrix_A[12210],matrix_B[10],mul_res1[12210]);
multi_7x28 multi_7x28_mod_12211(clk,rst,matrix_A[12211],matrix_B[11],mul_res1[12211]);
multi_7x28 multi_7x28_mod_12212(clk,rst,matrix_A[12212],matrix_B[12],mul_res1[12212]);
multi_7x28 multi_7x28_mod_12213(clk,rst,matrix_A[12213],matrix_B[13],mul_res1[12213]);
multi_7x28 multi_7x28_mod_12214(clk,rst,matrix_A[12214],matrix_B[14],mul_res1[12214]);
multi_7x28 multi_7x28_mod_12215(clk,rst,matrix_A[12215],matrix_B[15],mul_res1[12215]);
multi_7x28 multi_7x28_mod_12216(clk,rst,matrix_A[12216],matrix_B[16],mul_res1[12216]);
multi_7x28 multi_7x28_mod_12217(clk,rst,matrix_A[12217],matrix_B[17],mul_res1[12217]);
multi_7x28 multi_7x28_mod_12218(clk,rst,matrix_A[12218],matrix_B[18],mul_res1[12218]);
multi_7x28 multi_7x28_mod_12219(clk,rst,matrix_A[12219],matrix_B[19],mul_res1[12219]);
multi_7x28 multi_7x28_mod_12220(clk,rst,matrix_A[12220],matrix_B[20],mul_res1[12220]);
multi_7x28 multi_7x28_mod_12221(clk,rst,matrix_A[12221],matrix_B[21],mul_res1[12221]);
multi_7x28 multi_7x28_mod_12222(clk,rst,matrix_A[12222],matrix_B[22],mul_res1[12222]);
multi_7x28 multi_7x28_mod_12223(clk,rst,matrix_A[12223],matrix_B[23],mul_res1[12223]);
multi_7x28 multi_7x28_mod_12224(clk,rst,matrix_A[12224],matrix_B[24],mul_res1[12224]);
multi_7x28 multi_7x28_mod_12225(clk,rst,matrix_A[12225],matrix_B[25],mul_res1[12225]);
multi_7x28 multi_7x28_mod_12226(clk,rst,matrix_A[12226],matrix_B[26],mul_res1[12226]);
multi_7x28 multi_7x28_mod_12227(clk,rst,matrix_A[12227],matrix_B[27],mul_res1[12227]);
multi_7x28 multi_7x28_mod_12228(clk,rst,matrix_A[12228],matrix_B[28],mul_res1[12228]);
multi_7x28 multi_7x28_mod_12229(clk,rst,matrix_A[12229],matrix_B[29],mul_res1[12229]);
multi_7x28 multi_7x28_mod_12230(clk,rst,matrix_A[12230],matrix_B[30],mul_res1[12230]);
multi_7x28 multi_7x28_mod_12231(clk,rst,matrix_A[12231],matrix_B[31],mul_res1[12231]);
multi_7x28 multi_7x28_mod_12232(clk,rst,matrix_A[12232],matrix_B[32],mul_res1[12232]);
multi_7x28 multi_7x28_mod_12233(clk,rst,matrix_A[12233],matrix_B[33],mul_res1[12233]);
multi_7x28 multi_7x28_mod_12234(clk,rst,matrix_A[12234],matrix_B[34],mul_res1[12234]);
multi_7x28 multi_7x28_mod_12235(clk,rst,matrix_A[12235],matrix_B[35],mul_res1[12235]);
multi_7x28 multi_7x28_mod_12236(clk,rst,matrix_A[12236],matrix_B[36],mul_res1[12236]);
multi_7x28 multi_7x28_mod_12237(clk,rst,matrix_A[12237],matrix_B[37],mul_res1[12237]);
multi_7x28 multi_7x28_mod_12238(clk,rst,matrix_A[12238],matrix_B[38],mul_res1[12238]);
multi_7x28 multi_7x28_mod_12239(clk,rst,matrix_A[12239],matrix_B[39],mul_res1[12239]);
multi_7x28 multi_7x28_mod_12240(clk,rst,matrix_A[12240],matrix_B[40],mul_res1[12240]);
multi_7x28 multi_7x28_mod_12241(clk,rst,matrix_A[12241],matrix_B[41],mul_res1[12241]);
multi_7x28 multi_7x28_mod_12242(clk,rst,matrix_A[12242],matrix_B[42],mul_res1[12242]);
multi_7x28 multi_7x28_mod_12243(clk,rst,matrix_A[12243],matrix_B[43],mul_res1[12243]);
multi_7x28 multi_7x28_mod_12244(clk,rst,matrix_A[12244],matrix_B[44],mul_res1[12244]);
multi_7x28 multi_7x28_mod_12245(clk,rst,matrix_A[12245],matrix_B[45],mul_res1[12245]);
multi_7x28 multi_7x28_mod_12246(clk,rst,matrix_A[12246],matrix_B[46],mul_res1[12246]);
multi_7x28 multi_7x28_mod_12247(clk,rst,matrix_A[12247],matrix_B[47],mul_res1[12247]);
multi_7x28 multi_7x28_mod_12248(clk,rst,matrix_A[12248],matrix_B[48],mul_res1[12248]);
multi_7x28 multi_7x28_mod_12249(clk,rst,matrix_A[12249],matrix_B[49],mul_res1[12249]);
multi_7x28 multi_7x28_mod_12250(clk,rst,matrix_A[12250],matrix_B[50],mul_res1[12250]);
multi_7x28 multi_7x28_mod_12251(clk,rst,matrix_A[12251],matrix_B[51],mul_res1[12251]);
multi_7x28 multi_7x28_mod_12252(clk,rst,matrix_A[12252],matrix_B[52],mul_res1[12252]);
multi_7x28 multi_7x28_mod_12253(clk,rst,matrix_A[12253],matrix_B[53],mul_res1[12253]);
multi_7x28 multi_7x28_mod_12254(clk,rst,matrix_A[12254],matrix_B[54],mul_res1[12254]);
multi_7x28 multi_7x28_mod_12255(clk,rst,matrix_A[12255],matrix_B[55],mul_res1[12255]);
multi_7x28 multi_7x28_mod_12256(clk,rst,matrix_A[12256],matrix_B[56],mul_res1[12256]);
multi_7x28 multi_7x28_mod_12257(clk,rst,matrix_A[12257],matrix_B[57],mul_res1[12257]);
multi_7x28 multi_7x28_mod_12258(clk,rst,matrix_A[12258],matrix_B[58],mul_res1[12258]);
multi_7x28 multi_7x28_mod_12259(clk,rst,matrix_A[12259],matrix_B[59],mul_res1[12259]);
multi_7x28 multi_7x28_mod_12260(clk,rst,matrix_A[12260],matrix_B[60],mul_res1[12260]);
multi_7x28 multi_7x28_mod_12261(clk,rst,matrix_A[12261],matrix_B[61],mul_res1[12261]);
multi_7x28 multi_7x28_mod_12262(clk,rst,matrix_A[12262],matrix_B[62],mul_res1[12262]);
multi_7x28 multi_7x28_mod_12263(clk,rst,matrix_A[12263],matrix_B[63],mul_res1[12263]);
multi_7x28 multi_7x28_mod_12264(clk,rst,matrix_A[12264],matrix_B[64],mul_res1[12264]);
multi_7x28 multi_7x28_mod_12265(clk,rst,matrix_A[12265],matrix_B[65],mul_res1[12265]);
multi_7x28 multi_7x28_mod_12266(clk,rst,matrix_A[12266],matrix_B[66],mul_res1[12266]);
multi_7x28 multi_7x28_mod_12267(clk,rst,matrix_A[12267],matrix_B[67],mul_res1[12267]);
multi_7x28 multi_7x28_mod_12268(clk,rst,matrix_A[12268],matrix_B[68],mul_res1[12268]);
multi_7x28 multi_7x28_mod_12269(clk,rst,matrix_A[12269],matrix_B[69],mul_res1[12269]);
multi_7x28 multi_7x28_mod_12270(clk,rst,matrix_A[12270],matrix_B[70],mul_res1[12270]);
multi_7x28 multi_7x28_mod_12271(clk,rst,matrix_A[12271],matrix_B[71],mul_res1[12271]);
multi_7x28 multi_7x28_mod_12272(clk,rst,matrix_A[12272],matrix_B[72],mul_res1[12272]);
multi_7x28 multi_7x28_mod_12273(clk,rst,matrix_A[12273],matrix_B[73],mul_res1[12273]);
multi_7x28 multi_7x28_mod_12274(clk,rst,matrix_A[12274],matrix_B[74],mul_res1[12274]);
multi_7x28 multi_7x28_mod_12275(clk,rst,matrix_A[12275],matrix_B[75],mul_res1[12275]);
multi_7x28 multi_7x28_mod_12276(clk,rst,matrix_A[12276],matrix_B[76],mul_res1[12276]);
multi_7x28 multi_7x28_mod_12277(clk,rst,matrix_A[12277],matrix_B[77],mul_res1[12277]);
multi_7x28 multi_7x28_mod_12278(clk,rst,matrix_A[12278],matrix_B[78],mul_res1[12278]);
multi_7x28 multi_7x28_mod_12279(clk,rst,matrix_A[12279],matrix_B[79],mul_res1[12279]);
multi_7x28 multi_7x28_mod_12280(clk,rst,matrix_A[12280],matrix_B[80],mul_res1[12280]);
multi_7x28 multi_7x28_mod_12281(clk,rst,matrix_A[12281],matrix_B[81],mul_res1[12281]);
multi_7x28 multi_7x28_mod_12282(clk,rst,matrix_A[12282],matrix_B[82],mul_res1[12282]);
multi_7x28 multi_7x28_mod_12283(clk,rst,matrix_A[12283],matrix_B[83],mul_res1[12283]);
multi_7x28 multi_7x28_mod_12284(clk,rst,matrix_A[12284],matrix_B[84],mul_res1[12284]);
multi_7x28 multi_7x28_mod_12285(clk,rst,matrix_A[12285],matrix_B[85],mul_res1[12285]);
multi_7x28 multi_7x28_mod_12286(clk,rst,matrix_A[12286],matrix_B[86],mul_res1[12286]);
multi_7x28 multi_7x28_mod_12287(clk,rst,matrix_A[12287],matrix_B[87],mul_res1[12287]);
multi_7x28 multi_7x28_mod_12288(clk,rst,matrix_A[12288],matrix_B[88],mul_res1[12288]);
multi_7x28 multi_7x28_mod_12289(clk,rst,matrix_A[12289],matrix_B[89],mul_res1[12289]);
multi_7x28 multi_7x28_mod_12290(clk,rst,matrix_A[12290],matrix_B[90],mul_res1[12290]);
multi_7x28 multi_7x28_mod_12291(clk,rst,matrix_A[12291],matrix_B[91],mul_res1[12291]);
multi_7x28 multi_7x28_mod_12292(clk,rst,matrix_A[12292],matrix_B[92],mul_res1[12292]);
multi_7x28 multi_7x28_mod_12293(clk,rst,matrix_A[12293],matrix_B[93],mul_res1[12293]);
multi_7x28 multi_7x28_mod_12294(clk,rst,matrix_A[12294],matrix_B[94],mul_res1[12294]);
multi_7x28 multi_7x28_mod_12295(clk,rst,matrix_A[12295],matrix_B[95],mul_res1[12295]);
multi_7x28 multi_7x28_mod_12296(clk,rst,matrix_A[12296],matrix_B[96],mul_res1[12296]);
multi_7x28 multi_7x28_mod_12297(clk,rst,matrix_A[12297],matrix_B[97],mul_res1[12297]);
multi_7x28 multi_7x28_mod_12298(clk,rst,matrix_A[12298],matrix_B[98],mul_res1[12298]);
multi_7x28 multi_7x28_mod_12299(clk,rst,matrix_A[12299],matrix_B[99],mul_res1[12299]);
multi_7x28 multi_7x28_mod_12300(clk,rst,matrix_A[12300],matrix_B[100],mul_res1[12300]);
multi_7x28 multi_7x28_mod_12301(clk,rst,matrix_A[12301],matrix_B[101],mul_res1[12301]);
multi_7x28 multi_7x28_mod_12302(clk,rst,matrix_A[12302],matrix_B[102],mul_res1[12302]);
multi_7x28 multi_7x28_mod_12303(clk,rst,matrix_A[12303],matrix_B[103],mul_res1[12303]);
multi_7x28 multi_7x28_mod_12304(clk,rst,matrix_A[12304],matrix_B[104],mul_res1[12304]);
multi_7x28 multi_7x28_mod_12305(clk,rst,matrix_A[12305],matrix_B[105],mul_res1[12305]);
multi_7x28 multi_7x28_mod_12306(clk,rst,matrix_A[12306],matrix_B[106],mul_res1[12306]);
multi_7x28 multi_7x28_mod_12307(clk,rst,matrix_A[12307],matrix_B[107],mul_res1[12307]);
multi_7x28 multi_7x28_mod_12308(clk,rst,matrix_A[12308],matrix_B[108],mul_res1[12308]);
multi_7x28 multi_7x28_mod_12309(clk,rst,matrix_A[12309],matrix_B[109],mul_res1[12309]);
multi_7x28 multi_7x28_mod_12310(clk,rst,matrix_A[12310],matrix_B[110],mul_res1[12310]);
multi_7x28 multi_7x28_mod_12311(clk,rst,matrix_A[12311],matrix_B[111],mul_res1[12311]);
multi_7x28 multi_7x28_mod_12312(clk,rst,matrix_A[12312],matrix_B[112],mul_res1[12312]);
multi_7x28 multi_7x28_mod_12313(clk,rst,matrix_A[12313],matrix_B[113],mul_res1[12313]);
multi_7x28 multi_7x28_mod_12314(clk,rst,matrix_A[12314],matrix_B[114],mul_res1[12314]);
multi_7x28 multi_7x28_mod_12315(clk,rst,matrix_A[12315],matrix_B[115],mul_res1[12315]);
multi_7x28 multi_7x28_mod_12316(clk,rst,matrix_A[12316],matrix_B[116],mul_res1[12316]);
multi_7x28 multi_7x28_mod_12317(clk,rst,matrix_A[12317],matrix_B[117],mul_res1[12317]);
multi_7x28 multi_7x28_mod_12318(clk,rst,matrix_A[12318],matrix_B[118],mul_res1[12318]);
multi_7x28 multi_7x28_mod_12319(clk,rst,matrix_A[12319],matrix_B[119],mul_res1[12319]);
multi_7x28 multi_7x28_mod_12320(clk,rst,matrix_A[12320],matrix_B[120],mul_res1[12320]);
multi_7x28 multi_7x28_mod_12321(clk,rst,matrix_A[12321],matrix_B[121],mul_res1[12321]);
multi_7x28 multi_7x28_mod_12322(clk,rst,matrix_A[12322],matrix_B[122],mul_res1[12322]);
multi_7x28 multi_7x28_mod_12323(clk,rst,matrix_A[12323],matrix_B[123],mul_res1[12323]);
multi_7x28 multi_7x28_mod_12324(clk,rst,matrix_A[12324],matrix_B[124],mul_res1[12324]);
multi_7x28 multi_7x28_mod_12325(clk,rst,matrix_A[12325],matrix_B[125],mul_res1[12325]);
multi_7x28 multi_7x28_mod_12326(clk,rst,matrix_A[12326],matrix_B[126],mul_res1[12326]);
multi_7x28 multi_7x28_mod_12327(clk,rst,matrix_A[12327],matrix_B[127],mul_res1[12327]);
multi_7x28 multi_7x28_mod_12328(clk,rst,matrix_A[12328],matrix_B[128],mul_res1[12328]);
multi_7x28 multi_7x28_mod_12329(clk,rst,matrix_A[12329],matrix_B[129],mul_res1[12329]);
multi_7x28 multi_7x28_mod_12330(clk,rst,matrix_A[12330],matrix_B[130],mul_res1[12330]);
multi_7x28 multi_7x28_mod_12331(clk,rst,matrix_A[12331],matrix_B[131],mul_res1[12331]);
multi_7x28 multi_7x28_mod_12332(clk,rst,matrix_A[12332],matrix_B[132],mul_res1[12332]);
multi_7x28 multi_7x28_mod_12333(clk,rst,matrix_A[12333],matrix_B[133],mul_res1[12333]);
multi_7x28 multi_7x28_mod_12334(clk,rst,matrix_A[12334],matrix_B[134],mul_res1[12334]);
multi_7x28 multi_7x28_mod_12335(clk,rst,matrix_A[12335],matrix_B[135],mul_res1[12335]);
multi_7x28 multi_7x28_mod_12336(clk,rst,matrix_A[12336],matrix_B[136],mul_res1[12336]);
multi_7x28 multi_7x28_mod_12337(clk,rst,matrix_A[12337],matrix_B[137],mul_res1[12337]);
multi_7x28 multi_7x28_mod_12338(clk,rst,matrix_A[12338],matrix_B[138],mul_res1[12338]);
multi_7x28 multi_7x28_mod_12339(clk,rst,matrix_A[12339],matrix_B[139],mul_res1[12339]);
multi_7x28 multi_7x28_mod_12340(clk,rst,matrix_A[12340],matrix_B[140],mul_res1[12340]);
multi_7x28 multi_7x28_mod_12341(clk,rst,matrix_A[12341],matrix_B[141],mul_res1[12341]);
multi_7x28 multi_7x28_mod_12342(clk,rst,matrix_A[12342],matrix_B[142],mul_res1[12342]);
multi_7x28 multi_7x28_mod_12343(clk,rst,matrix_A[12343],matrix_B[143],mul_res1[12343]);
multi_7x28 multi_7x28_mod_12344(clk,rst,matrix_A[12344],matrix_B[144],mul_res1[12344]);
multi_7x28 multi_7x28_mod_12345(clk,rst,matrix_A[12345],matrix_B[145],mul_res1[12345]);
multi_7x28 multi_7x28_mod_12346(clk,rst,matrix_A[12346],matrix_B[146],mul_res1[12346]);
multi_7x28 multi_7x28_mod_12347(clk,rst,matrix_A[12347],matrix_B[147],mul_res1[12347]);
multi_7x28 multi_7x28_mod_12348(clk,rst,matrix_A[12348],matrix_B[148],mul_res1[12348]);
multi_7x28 multi_7x28_mod_12349(clk,rst,matrix_A[12349],matrix_B[149],mul_res1[12349]);
multi_7x28 multi_7x28_mod_12350(clk,rst,matrix_A[12350],matrix_B[150],mul_res1[12350]);
multi_7x28 multi_7x28_mod_12351(clk,rst,matrix_A[12351],matrix_B[151],mul_res1[12351]);
multi_7x28 multi_7x28_mod_12352(clk,rst,matrix_A[12352],matrix_B[152],mul_res1[12352]);
multi_7x28 multi_7x28_mod_12353(clk,rst,matrix_A[12353],matrix_B[153],mul_res1[12353]);
multi_7x28 multi_7x28_mod_12354(clk,rst,matrix_A[12354],matrix_B[154],mul_res1[12354]);
multi_7x28 multi_7x28_mod_12355(clk,rst,matrix_A[12355],matrix_B[155],mul_res1[12355]);
multi_7x28 multi_7x28_mod_12356(clk,rst,matrix_A[12356],matrix_B[156],mul_res1[12356]);
multi_7x28 multi_7x28_mod_12357(clk,rst,matrix_A[12357],matrix_B[157],mul_res1[12357]);
multi_7x28 multi_7x28_mod_12358(clk,rst,matrix_A[12358],matrix_B[158],mul_res1[12358]);
multi_7x28 multi_7x28_mod_12359(clk,rst,matrix_A[12359],matrix_B[159],mul_res1[12359]);
multi_7x28 multi_7x28_mod_12360(clk,rst,matrix_A[12360],matrix_B[160],mul_res1[12360]);
multi_7x28 multi_7x28_mod_12361(clk,rst,matrix_A[12361],matrix_B[161],mul_res1[12361]);
multi_7x28 multi_7x28_mod_12362(clk,rst,matrix_A[12362],matrix_B[162],mul_res1[12362]);
multi_7x28 multi_7x28_mod_12363(clk,rst,matrix_A[12363],matrix_B[163],mul_res1[12363]);
multi_7x28 multi_7x28_mod_12364(clk,rst,matrix_A[12364],matrix_B[164],mul_res1[12364]);
multi_7x28 multi_7x28_mod_12365(clk,rst,matrix_A[12365],matrix_B[165],mul_res1[12365]);
multi_7x28 multi_7x28_mod_12366(clk,rst,matrix_A[12366],matrix_B[166],mul_res1[12366]);
multi_7x28 multi_7x28_mod_12367(clk,rst,matrix_A[12367],matrix_B[167],mul_res1[12367]);
multi_7x28 multi_7x28_mod_12368(clk,rst,matrix_A[12368],matrix_B[168],mul_res1[12368]);
multi_7x28 multi_7x28_mod_12369(clk,rst,matrix_A[12369],matrix_B[169],mul_res1[12369]);
multi_7x28 multi_7x28_mod_12370(clk,rst,matrix_A[12370],matrix_B[170],mul_res1[12370]);
multi_7x28 multi_7x28_mod_12371(clk,rst,matrix_A[12371],matrix_B[171],mul_res1[12371]);
multi_7x28 multi_7x28_mod_12372(clk,rst,matrix_A[12372],matrix_B[172],mul_res1[12372]);
multi_7x28 multi_7x28_mod_12373(clk,rst,matrix_A[12373],matrix_B[173],mul_res1[12373]);
multi_7x28 multi_7x28_mod_12374(clk,rst,matrix_A[12374],matrix_B[174],mul_res1[12374]);
multi_7x28 multi_7x28_mod_12375(clk,rst,matrix_A[12375],matrix_B[175],mul_res1[12375]);
multi_7x28 multi_7x28_mod_12376(clk,rst,matrix_A[12376],matrix_B[176],mul_res1[12376]);
multi_7x28 multi_7x28_mod_12377(clk,rst,matrix_A[12377],matrix_B[177],mul_res1[12377]);
multi_7x28 multi_7x28_mod_12378(clk,rst,matrix_A[12378],matrix_B[178],mul_res1[12378]);
multi_7x28 multi_7x28_mod_12379(clk,rst,matrix_A[12379],matrix_B[179],mul_res1[12379]);
multi_7x28 multi_7x28_mod_12380(clk,rst,matrix_A[12380],matrix_B[180],mul_res1[12380]);
multi_7x28 multi_7x28_mod_12381(clk,rst,matrix_A[12381],matrix_B[181],mul_res1[12381]);
multi_7x28 multi_7x28_mod_12382(clk,rst,matrix_A[12382],matrix_B[182],mul_res1[12382]);
multi_7x28 multi_7x28_mod_12383(clk,rst,matrix_A[12383],matrix_B[183],mul_res1[12383]);
multi_7x28 multi_7x28_mod_12384(clk,rst,matrix_A[12384],matrix_B[184],mul_res1[12384]);
multi_7x28 multi_7x28_mod_12385(clk,rst,matrix_A[12385],matrix_B[185],mul_res1[12385]);
multi_7x28 multi_7x28_mod_12386(clk,rst,matrix_A[12386],matrix_B[186],mul_res1[12386]);
multi_7x28 multi_7x28_mod_12387(clk,rst,matrix_A[12387],matrix_B[187],mul_res1[12387]);
multi_7x28 multi_7x28_mod_12388(clk,rst,matrix_A[12388],matrix_B[188],mul_res1[12388]);
multi_7x28 multi_7x28_mod_12389(clk,rst,matrix_A[12389],matrix_B[189],mul_res1[12389]);
multi_7x28 multi_7x28_mod_12390(clk,rst,matrix_A[12390],matrix_B[190],mul_res1[12390]);
multi_7x28 multi_7x28_mod_12391(clk,rst,matrix_A[12391],matrix_B[191],mul_res1[12391]);
multi_7x28 multi_7x28_mod_12392(clk,rst,matrix_A[12392],matrix_B[192],mul_res1[12392]);
multi_7x28 multi_7x28_mod_12393(clk,rst,matrix_A[12393],matrix_B[193],mul_res1[12393]);
multi_7x28 multi_7x28_mod_12394(clk,rst,matrix_A[12394],matrix_B[194],mul_res1[12394]);
multi_7x28 multi_7x28_mod_12395(clk,rst,matrix_A[12395],matrix_B[195],mul_res1[12395]);
multi_7x28 multi_7x28_mod_12396(clk,rst,matrix_A[12396],matrix_B[196],mul_res1[12396]);
multi_7x28 multi_7x28_mod_12397(clk,rst,matrix_A[12397],matrix_B[197],mul_res1[12397]);
multi_7x28 multi_7x28_mod_12398(clk,rst,matrix_A[12398],matrix_B[198],mul_res1[12398]);
multi_7x28 multi_7x28_mod_12399(clk,rst,matrix_A[12399],matrix_B[199],mul_res1[12399]);
multi_7x28 multi_7x28_mod_12400(clk,rst,matrix_A[12400],matrix_B[0],mul_res1[12400]);
multi_7x28 multi_7x28_mod_12401(clk,rst,matrix_A[12401],matrix_B[1],mul_res1[12401]);
multi_7x28 multi_7x28_mod_12402(clk,rst,matrix_A[12402],matrix_B[2],mul_res1[12402]);
multi_7x28 multi_7x28_mod_12403(clk,rst,matrix_A[12403],matrix_B[3],mul_res1[12403]);
multi_7x28 multi_7x28_mod_12404(clk,rst,matrix_A[12404],matrix_B[4],mul_res1[12404]);
multi_7x28 multi_7x28_mod_12405(clk,rst,matrix_A[12405],matrix_B[5],mul_res1[12405]);
multi_7x28 multi_7x28_mod_12406(clk,rst,matrix_A[12406],matrix_B[6],mul_res1[12406]);
multi_7x28 multi_7x28_mod_12407(clk,rst,matrix_A[12407],matrix_B[7],mul_res1[12407]);
multi_7x28 multi_7x28_mod_12408(clk,rst,matrix_A[12408],matrix_B[8],mul_res1[12408]);
multi_7x28 multi_7x28_mod_12409(clk,rst,matrix_A[12409],matrix_B[9],mul_res1[12409]);
multi_7x28 multi_7x28_mod_12410(clk,rst,matrix_A[12410],matrix_B[10],mul_res1[12410]);
multi_7x28 multi_7x28_mod_12411(clk,rst,matrix_A[12411],matrix_B[11],mul_res1[12411]);
multi_7x28 multi_7x28_mod_12412(clk,rst,matrix_A[12412],matrix_B[12],mul_res1[12412]);
multi_7x28 multi_7x28_mod_12413(clk,rst,matrix_A[12413],matrix_B[13],mul_res1[12413]);
multi_7x28 multi_7x28_mod_12414(clk,rst,matrix_A[12414],matrix_B[14],mul_res1[12414]);
multi_7x28 multi_7x28_mod_12415(clk,rst,matrix_A[12415],matrix_B[15],mul_res1[12415]);
multi_7x28 multi_7x28_mod_12416(clk,rst,matrix_A[12416],matrix_B[16],mul_res1[12416]);
multi_7x28 multi_7x28_mod_12417(clk,rst,matrix_A[12417],matrix_B[17],mul_res1[12417]);
multi_7x28 multi_7x28_mod_12418(clk,rst,matrix_A[12418],matrix_B[18],mul_res1[12418]);
multi_7x28 multi_7x28_mod_12419(clk,rst,matrix_A[12419],matrix_B[19],mul_res1[12419]);
multi_7x28 multi_7x28_mod_12420(clk,rst,matrix_A[12420],matrix_B[20],mul_res1[12420]);
multi_7x28 multi_7x28_mod_12421(clk,rst,matrix_A[12421],matrix_B[21],mul_res1[12421]);
multi_7x28 multi_7x28_mod_12422(clk,rst,matrix_A[12422],matrix_B[22],mul_res1[12422]);
multi_7x28 multi_7x28_mod_12423(clk,rst,matrix_A[12423],matrix_B[23],mul_res1[12423]);
multi_7x28 multi_7x28_mod_12424(clk,rst,matrix_A[12424],matrix_B[24],mul_res1[12424]);
multi_7x28 multi_7x28_mod_12425(clk,rst,matrix_A[12425],matrix_B[25],mul_res1[12425]);
multi_7x28 multi_7x28_mod_12426(clk,rst,matrix_A[12426],matrix_B[26],mul_res1[12426]);
multi_7x28 multi_7x28_mod_12427(clk,rst,matrix_A[12427],matrix_B[27],mul_res1[12427]);
multi_7x28 multi_7x28_mod_12428(clk,rst,matrix_A[12428],matrix_B[28],mul_res1[12428]);
multi_7x28 multi_7x28_mod_12429(clk,rst,matrix_A[12429],matrix_B[29],mul_res1[12429]);
multi_7x28 multi_7x28_mod_12430(clk,rst,matrix_A[12430],matrix_B[30],mul_res1[12430]);
multi_7x28 multi_7x28_mod_12431(clk,rst,matrix_A[12431],matrix_B[31],mul_res1[12431]);
multi_7x28 multi_7x28_mod_12432(clk,rst,matrix_A[12432],matrix_B[32],mul_res1[12432]);
multi_7x28 multi_7x28_mod_12433(clk,rst,matrix_A[12433],matrix_B[33],mul_res1[12433]);
multi_7x28 multi_7x28_mod_12434(clk,rst,matrix_A[12434],matrix_B[34],mul_res1[12434]);
multi_7x28 multi_7x28_mod_12435(clk,rst,matrix_A[12435],matrix_B[35],mul_res1[12435]);
multi_7x28 multi_7x28_mod_12436(clk,rst,matrix_A[12436],matrix_B[36],mul_res1[12436]);
multi_7x28 multi_7x28_mod_12437(clk,rst,matrix_A[12437],matrix_B[37],mul_res1[12437]);
multi_7x28 multi_7x28_mod_12438(clk,rst,matrix_A[12438],matrix_B[38],mul_res1[12438]);
multi_7x28 multi_7x28_mod_12439(clk,rst,matrix_A[12439],matrix_B[39],mul_res1[12439]);
multi_7x28 multi_7x28_mod_12440(clk,rst,matrix_A[12440],matrix_B[40],mul_res1[12440]);
multi_7x28 multi_7x28_mod_12441(clk,rst,matrix_A[12441],matrix_B[41],mul_res1[12441]);
multi_7x28 multi_7x28_mod_12442(clk,rst,matrix_A[12442],matrix_B[42],mul_res1[12442]);
multi_7x28 multi_7x28_mod_12443(clk,rst,matrix_A[12443],matrix_B[43],mul_res1[12443]);
multi_7x28 multi_7x28_mod_12444(clk,rst,matrix_A[12444],matrix_B[44],mul_res1[12444]);
multi_7x28 multi_7x28_mod_12445(clk,rst,matrix_A[12445],matrix_B[45],mul_res1[12445]);
multi_7x28 multi_7x28_mod_12446(clk,rst,matrix_A[12446],matrix_B[46],mul_res1[12446]);
multi_7x28 multi_7x28_mod_12447(clk,rst,matrix_A[12447],matrix_B[47],mul_res1[12447]);
multi_7x28 multi_7x28_mod_12448(clk,rst,matrix_A[12448],matrix_B[48],mul_res1[12448]);
multi_7x28 multi_7x28_mod_12449(clk,rst,matrix_A[12449],matrix_B[49],mul_res1[12449]);
multi_7x28 multi_7x28_mod_12450(clk,rst,matrix_A[12450],matrix_B[50],mul_res1[12450]);
multi_7x28 multi_7x28_mod_12451(clk,rst,matrix_A[12451],matrix_B[51],mul_res1[12451]);
multi_7x28 multi_7x28_mod_12452(clk,rst,matrix_A[12452],matrix_B[52],mul_res1[12452]);
multi_7x28 multi_7x28_mod_12453(clk,rst,matrix_A[12453],matrix_B[53],mul_res1[12453]);
multi_7x28 multi_7x28_mod_12454(clk,rst,matrix_A[12454],matrix_B[54],mul_res1[12454]);
multi_7x28 multi_7x28_mod_12455(clk,rst,matrix_A[12455],matrix_B[55],mul_res1[12455]);
multi_7x28 multi_7x28_mod_12456(clk,rst,matrix_A[12456],matrix_B[56],mul_res1[12456]);
multi_7x28 multi_7x28_mod_12457(clk,rst,matrix_A[12457],matrix_B[57],mul_res1[12457]);
multi_7x28 multi_7x28_mod_12458(clk,rst,matrix_A[12458],matrix_B[58],mul_res1[12458]);
multi_7x28 multi_7x28_mod_12459(clk,rst,matrix_A[12459],matrix_B[59],mul_res1[12459]);
multi_7x28 multi_7x28_mod_12460(clk,rst,matrix_A[12460],matrix_B[60],mul_res1[12460]);
multi_7x28 multi_7x28_mod_12461(clk,rst,matrix_A[12461],matrix_B[61],mul_res1[12461]);
multi_7x28 multi_7x28_mod_12462(clk,rst,matrix_A[12462],matrix_B[62],mul_res1[12462]);
multi_7x28 multi_7x28_mod_12463(clk,rst,matrix_A[12463],matrix_B[63],mul_res1[12463]);
multi_7x28 multi_7x28_mod_12464(clk,rst,matrix_A[12464],matrix_B[64],mul_res1[12464]);
multi_7x28 multi_7x28_mod_12465(clk,rst,matrix_A[12465],matrix_B[65],mul_res1[12465]);
multi_7x28 multi_7x28_mod_12466(clk,rst,matrix_A[12466],matrix_B[66],mul_res1[12466]);
multi_7x28 multi_7x28_mod_12467(clk,rst,matrix_A[12467],matrix_B[67],mul_res1[12467]);
multi_7x28 multi_7x28_mod_12468(clk,rst,matrix_A[12468],matrix_B[68],mul_res1[12468]);
multi_7x28 multi_7x28_mod_12469(clk,rst,matrix_A[12469],matrix_B[69],mul_res1[12469]);
multi_7x28 multi_7x28_mod_12470(clk,rst,matrix_A[12470],matrix_B[70],mul_res1[12470]);
multi_7x28 multi_7x28_mod_12471(clk,rst,matrix_A[12471],matrix_B[71],mul_res1[12471]);
multi_7x28 multi_7x28_mod_12472(clk,rst,matrix_A[12472],matrix_B[72],mul_res1[12472]);
multi_7x28 multi_7x28_mod_12473(clk,rst,matrix_A[12473],matrix_B[73],mul_res1[12473]);
multi_7x28 multi_7x28_mod_12474(clk,rst,matrix_A[12474],matrix_B[74],mul_res1[12474]);
multi_7x28 multi_7x28_mod_12475(clk,rst,matrix_A[12475],matrix_B[75],mul_res1[12475]);
multi_7x28 multi_7x28_mod_12476(clk,rst,matrix_A[12476],matrix_B[76],mul_res1[12476]);
multi_7x28 multi_7x28_mod_12477(clk,rst,matrix_A[12477],matrix_B[77],mul_res1[12477]);
multi_7x28 multi_7x28_mod_12478(clk,rst,matrix_A[12478],matrix_B[78],mul_res1[12478]);
multi_7x28 multi_7x28_mod_12479(clk,rst,matrix_A[12479],matrix_B[79],mul_res1[12479]);
multi_7x28 multi_7x28_mod_12480(clk,rst,matrix_A[12480],matrix_B[80],mul_res1[12480]);
multi_7x28 multi_7x28_mod_12481(clk,rst,matrix_A[12481],matrix_B[81],mul_res1[12481]);
multi_7x28 multi_7x28_mod_12482(clk,rst,matrix_A[12482],matrix_B[82],mul_res1[12482]);
multi_7x28 multi_7x28_mod_12483(clk,rst,matrix_A[12483],matrix_B[83],mul_res1[12483]);
multi_7x28 multi_7x28_mod_12484(clk,rst,matrix_A[12484],matrix_B[84],mul_res1[12484]);
multi_7x28 multi_7x28_mod_12485(clk,rst,matrix_A[12485],matrix_B[85],mul_res1[12485]);
multi_7x28 multi_7x28_mod_12486(clk,rst,matrix_A[12486],matrix_B[86],mul_res1[12486]);
multi_7x28 multi_7x28_mod_12487(clk,rst,matrix_A[12487],matrix_B[87],mul_res1[12487]);
multi_7x28 multi_7x28_mod_12488(clk,rst,matrix_A[12488],matrix_B[88],mul_res1[12488]);
multi_7x28 multi_7x28_mod_12489(clk,rst,matrix_A[12489],matrix_B[89],mul_res1[12489]);
multi_7x28 multi_7x28_mod_12490(clk,rst,matrix_A[12490],matrix_B[90],mul_res1[12490]);
multi_7x28 multi_7x28_mod_12491(clk,rst,matrix_A[12491],matrix_B[91],mul_res1[12491]);
multi_7x28 multi_7x28_mod_12492(clk,rst,matrix_A[12492],matrix_B[92],mul_res1[12492]);
multi_7x28 multi_7x28_mod_12493(clk,rst,matrix_A[12493],matrix_B[93],mul_res1[12493]);
multi_7x28 multi_7x28_mod_12494(clk,rst,matrix_A[12494],matrix_B[94],mul_res1[12494]);
multi_7x28 multi_7x28_mod_12495(clk,rst,matrix_A[12495],matrix_B[95],mul_res1[12495]);
multi_7x28 multi_7x28_mod_12496(clk,rst,matrix_A[12496],matrix_B[96],mul_res1[12496]);
multi_7x28 multi_7x28_mod_12497(clk,rst,matrix_A[12497],matrix_B[97],mul_res1[12497]);
multi_7x28 multi_7x28_mod_12498(clk,rst,matrix_A[12498],matrix_B[98],mul_res1[12498]);
multi_7x28 multi_7x28_mod_12499(clk,rst,matrix_A[12499],matrix_B[99],mul_res1[12499]);
multi_7x28 multi_7x28_mod_12500(clk,rst,matrix_A[12500],matrix_B[100],mul_res1[12500]);
multi_7x28 multi_7x28_mod_12501(clk,rst,matrix_A[12501],matrix_B[101],mul_res1[12501]);
multi_7x28 multi_7x28_mod_12502(clk,rst,matrix_A[12502],matrix_B[102],mul_res1[12502]);
multi_7x28 multi_7x28_mod_12503(clk,rst,matrix_A[12503],matrix_B[103],mul_res1[12503]);
multi_7x28 multi_7x28_mod_12504(clk,rst,matrix_A[12504],matrix_B[104],mul_res1[12504]);
multi_7x28 multi_7x28_mod_12505(clk,rst,matrix_A[12505],matrix_B[105],mul_res1[12505]);
multi_7x28 multi_7x28_mod_12506(clk,rst,matrix_A[12506],matrix_B[106],mul_res1[12506]);
multi_7x28 multi_7x28_mod_12507(clk,rst,matrix_A[12507],matrix_B[107],mul_res1[12507]);
multi_7x28 multi_7x28_mod_12508(clk,rst,matrix_A[12508],matrix_B[108],mul_res1[12508]);
multi_7x28 multi_7x28_mod_12509(clk,rst,matrix_A[12509],matrix_B[109],mul_res1[12509]);
multi_7x28 multi_7x28_mod_12510(clk,rst,matrix_A[12510],matrix_B[110],mul_res1[12510]);
multi_7x28 multi_7x28_mod_12511(clk,rst,matrix_A[12511],matrix_B[111],mul_res1[12511]);
multi_7x28 multi_7x28_mod_12512(clk,rst,matrix_A[12512],matrix_B[112],mul_res1[12512]);
multi_7x28 multi_7x28_mod_12513(clk,rst,matrix_A[12513],matrix_B[113],mul_res1[12513]);
multi_7x28 multi_7x28_mod_12514(clk,rst,matrix_A[12514],matrix_B[114],mul_res1[12514]);
multi_7x28 multi_7x28_mod_12515(clk,rst,matrix_A[12515],matrix_B[115],mul_res1[12515]);
multi_7x28 multi_7x28_mod_12516(clk,rst,matrix_A[12516],matrix_B[116],mul_res1[12516]);
multi_7x28 multi_7x28_mod_12517(clk,rst,matrix_A[12517],matrix_B[117],mul_res1[12517]);
multi_7x28 multi_7x28_mod_12518(clk,rst,matrix_A[12518],matrix_B[118],mul_res1[12518]);
multi_7x28 multi_7x28_mod_12519(clk,rst,matrix_A[12519],matrix_B[119],mul_res1[12519]);
multi_7x28 multi_7x28_mod_12520(clk,rst,matrix_A[12520],matrix_B[120],mul_res1[12520]);
multi_7x28 multi_7x28_mod_12521(clk,rst,matrix_A[12521],matrix_B[121],mul_res1[12521]);
multi_7x28 multi_7x28_mod_12522(clk,rst,matrix_A[12522],matrix_B[122],mul_res1[12522]);
multi_7x28 multi_7x28_mod_12523(clk,rst,matrix_A[12523],matrix_B[123],mul_res1[12523]);
multi_7x28 multi_7x28_mod_12524(clk,rst,matrix_A[12524],matrix_B[124],mul_res1[12524]);
multi_7x28 multi_7x28_mod_12525(clk,rst,matrix_A[12525],matrix_B[125],mul_res1[12525]);
multi_7x28 multi_7x28_mod_12526(clk,rst,matrix_A[12526],matrix_B[126],mul_res1[12526]);
multi_7x28 multi_7x28_mod_12527(clk,rst,matrix_A[12527],matrix_B[127],mul_res1[12527]);
multi_7x28 multi_7x28_mod_12528(clk,rst,matrix_A[12528],matrix_B[128],mul_res1[12528]);
multi_7x28 multi_7x28_mod_12529(clk,rst,matrix_A[12529],matrix_B[129],mul_res1[12529]);
multi_7x28 multi_7x28_mod_12530(clk,rst,matrix_A[12530],matrix_B[130],mul_res1[12530]);
multi_7x28 multi_7x28_mod_12531(clk,rst,matrix_A[12531],matrix_B[131],mul_res1[12531]);
multi_7x28 multi_7x28_mod_12532(clk,rst,matrix_A[12532],matrix_B[132],mul_res1[12532]);
multi_7x28 multi_7x28_mod_12533(clk,rst,matrix_A[12533],matrix_B[133],mul_res1[12533]);
multi_7x28 multi_7x28_mod_12534(clk,rst,matrix_A[12534],matrix_B[134],mul_res1[12534]);
multi_7x28 multi_7x28_mod_12535(clk,rst,matrix_A[12535],matrix_B[135],mul_res1[12535]);
multi_7x28 multi_7x28_mod_12536(clk,rst,matrix_A[12536],matrix_B[136],mul_res1[12536]);
multi_7x28 multi_7x28_mod_12537(clk,rst,matrix_A[12537],matrix_B[137],mul_res1[12537]);
multi_7x28 multi_7x28_mod_12538(clk,rst,matrix_A[12538],matrix_B[138],mul_res1[12538]);
multi_7x28 multi_7x28_mod_12539(clk,rst,matrix_A[12539],matrix_B[139],mul_res1[12539]);
multi_7x28 multi_7x28_mod_12540(clk,rst,matrix_A[12540],matrix_B[140],mul_res1[12540]);
multi_7x28 multi_7x28_mod_12541(clk,rst,matrix_A[12541],matrix_B[141],mul_res1[12541]);
multi_7x28 multi_7x28_mod_12542(clk,rst,matrix_A[12542],matrix_B[142],mul_res1[12542]);
multi_7x28 multi_7x28_mod_12543(clk,rst,matrix_A[12543],matrix_B[143],mul_res1[12543]);
multi_7x28 multi_7x28_mod_12544(clk,rst,matrix_A[12544],matrix_B[144],mul_res1[12544]);
multi_7x28 multi_7x28_mod_12545(clk,rst,matrix_A[12545],matrix_B[145],mul_res1[12545]);
multi_7x28 multi_7x28_mod_12546(clk,rst,matrix_A[12546],matrix_B[146],mul_res1[12546]);
multi_7x28 multi_7x28_mod_12547(clk,rst,matrix_A[12547],matrix_B[147],mul_res1[12547]);
multi_7x28 multi_7x28_mod_12548(clk,rst,matrix_A[12548],matrix_B[148],mul_res1[12548]);
multi_7x28 multi_7x28_mod_12549(clk,rst,matrix_A[12549],matrix_B[149],mul_res1[12549]);
multi_7x28 multi_7x28_mod_12550(clk,rst,matrix_A[12550],matrix_B[150],mul_res1[12550]);
multi_7x28 multi_7x28_mod_12551(clk,rst,matrix_A[12551],matrix_B[151],mul_res1[12551]);
multi_7x28 multi_7x28_mod_12552(clk,rst,matrix_A[12552],matrix_B[152],mul_res1[12552]);
multi_7x28 multi_7x28_mod_12553(clk,rst,matrix_A[12553],matrix_B[153],mul_res1[12553]);
multi_7x28 multi_7x28_mod_12554(clk,rst,matrix_A[12554],matrix_B[154],mul_res1[12554]);
multi_7x28 multi_7x28_mod_12555(clk,rst,matrix_A[12555],matrix_B[155],mul_res1[12555]);
multi_7x28 multi_7x28_mod_12556(clk,rst,matrix_A[12556],matrix_B[156],mul_res1[12556]);
multi_7x28 multi_7x28_mod_12557(clk,rst,matrix_A[12557],matrix_B[157],mul_res1[12557]);
multi_7x28 multi_7x28_mod_12558(clk,rst,matrix_A[12558],matrix_B[158],mul_res1[12558]);
multi_7x28 multi_7x28_mod_12559(clk,rst,matrix_A[12559],matrix_B[159],mul_res1[12559]);
multi_7x28 multi_7x28_mod_12560(clk,rst,matrix_A[12560],matrix_B[160],mul_res1[12560]);
multi_7x28 multi_7x28_mod_12561(clk,rst,matrix_A[12561],matrix_B[161],mul_res1[12561]);
multi_7x28 multi_7x28_mod_12562(clk,rst,matrix_A[12562],matrix_B[162],mul_res1[12562]);
multi_7x28 multi_7x28_mod_12563(clk,rst,matrix_A[12563],matrix_B[163],mul_res1[12563]);
multi_7x28 multi_7x28_mod_12564(clk,rst,matrix_A[12564],matrix_B[164],mul_res1[12564]);
multi_7x28 multi_7x28_mod_12565(clk,rst,matrix_A[12565],matrix_B[165],mul_res1[12565]);
multi_7x28 multi_7x28_mod_12566(clk,rst,matrix_A[12566],matrix_B[166],mul_res1[12566]);
multi_7x28 multi_7x28_mod_12567(clk,rst,matrix_A[12567],matrix_B[167],mul_res1[12567]);
multi_7x28 multi_7x28_mod_12568(clk,rst,matrix_A[12568],matrix_B[168],mul_res1[12568]);
multi_7x28 multi_7x28_mod_12569(clk,rst,matrix_A[12569],matrix_B[169],mul_res1[12569]);
multi_7x28 multi_7x28_mod_12570(clk,rst,matrix_A[12570],matrix_B[170],mul_res1[12570]);
multi_7x28 multi_7x28_mod_12571(clk,rst,matrix_A[12571],matrix_B[171],mul_res1[12571]);
multi_7x28 multi_7x28_mod_12572(clk,rst,matrix_A[12572],matrix_B[172],mul_res1[12572]);
multi_7x28 multi_7x28_mod_12573(clk,rst,matrix_A[12573],matrix_B[173],mul_res1[12573]);
multi_7x28 multi_7x28_mod_12574(clk,rst,matrix_A[12574],matrix_B[174],mul_res1[12574]);
multi_7x28 multi_7x28_mod_12575(clk,rst,matrix_A[12575],matrix_B[175],mul_res1[12575]);
multi_7x28 multi_7x28_mod_12576(clk,rst,matrix_A[12576],matrix_B[176],mul_res1[12576]);
multi_7x28 multi_7x28_mod_12577(clk,rst,matrix_A[12577],matrix_B[177],mul_res1[12577]);
multi_7x28 multi_7x28_mod_12578(clk,rst,matrix_A[12578],matrix_B[178],mul_res1[12578]);
multi_7x28 multi_7x28_mod_12579(clk,rst,matrix_A[12579],matrix_B[179],mul_res1[12579]);
multi_7x28 multi_7x28_mod_12580(clk,rst,matrix_A[12580],matrix_B[180],mul_res1[12580]);
multi_7x28 multi_7x28_mod_12581(clk,rst,matrix_A[12581],matrix_B[181],mul_res1[12581]);
multi_7x28 multi_7x28_mod_12582(clk,rst,matrix_A[12582],matrix_B[182],mul_res1[12582]);
multi_7x28 multi_7x28_mod_12583(clk,rst,matrix_A[12583],matrix_B[183],mul_res1[12583]);
multi_7x28 multi_7x28_mod_12584(clk,rst,matrix_A[12584],matrix_B[184],mul_res1[12584]);
multi_7x28 multi_7x28_mod_12585(clk,rst,matrix_A[12585],matrix_B[185],mul_res1[12585]);
multi_7x28 multi_7x28_mod_12586(clk,rst,matrix_A[12586],matrix_B[186],mul_res1[12586]);
multi_7x28 multi_7x28_mod_12587(clk,rst,matrix_A[12587],matrix_B[187],mul_res1[12587]);
multi_7x28 multi_7x28_mod_12588(clk,rst,matrix_A[12588],matrix_B[188],mul_res1[12588]);
multi_7x28 multi_7x28_mod_12589(clk,rst,matrix_A[12589],matrix_B[189],mul_res1[12589]);
multi_7x28 multi_7x28_mod_12590(clk,rst,matrix_A[12590],matrix_B[190],mul_res1[12590]);
multi_7x28 multi_7x28_mod_12591(clk,rst,matrix_A[12591],matrix_B[191],mul_res1[12591]);
multi_7x28 multi_7x28_mod_12592(clk,rst,matrix_A[12592],matrix_B[192],mul_res1[12592]);
multi_7x28 multi_7x28_mod_12593(clk,rst,matrix_A[12593],matrix_B[193],mul_res1[12593]);
multi_7x28 multi_7x28_mod_12594(clk,rst,matrix_A[12594],matrix_B[194],mul_res1[12594]);
multi_7x28 multi_7x28_mod_12595(clk,rst,matrix_A[12595],matrix_B[195],mul_res1[12595]);
multi_7x28 multi_7x28_mod_12596(clk,rst,matrix_A[12596],matrix_B[196],mul_res1[12596]);
multi_7x28 multi_7x28_mod_12597(clk,rst,matrix_A[12597],matrix_B[197],mul_res1[12597]);
multi_7x28 multi_7x28_mod_12598(clk,rst,matrix_A[12598],matrix_B[198],mul_res1[12598]);
multi_7x28 multi_7x28_mod_12599(clk,rst,matrix_A[12599],matrix_B[199],mul_res1[12599]);
multi_7x28 multi_7x28_mod_12600(clk,rst,matrix_A[12600],matrix_B[0],mul_res1[12600]);
multi_7x28 multi_7x28_mod_12601(clk,rst,matrix_A[12601],matrix_B[1],mul_res1[12601]);
multi_7x28 multi_7x28_mod_12602(clk,rst,matrix_A[12602],matrix_B[2],mul_res1[12602]);
multi_7x28 multi_7x28_mod_12603(clk,rst,matrix_A[12603],matrix_B[3],mul_res1[12603]);
multi_7x28 multi_7x28_mod_12604(clk,rst,matrix_A[12604],matrix_B[4],mul_res1[12604]);
multi_7x28 multi_7x28_mod_12605(clk,rst,matrix_A[12605],matrix_B[5],mul_res1[12605]);
multi_7x28 multi_7x28_mod_12606(clk,rst,matrix_A[12606],matrix_B[6],mul_res1[12606]);
multi_7x28 multi_7x28_mod_12607(clk,rst,matrix_A[12607],matrix_B[7],mul_res1[12607]);
multi_7x28 multi_7x28_mod_12608(clk,rst,matrix_A[12608],matrix_B[8],mul_res1[12608]);
multi_7x28 multi_7x28_mod_12609(clk,rst,matrix_A[12609],matrix_B[9],mul_res1[12609]);
multi_7x28 multi_7x28_mod_12610(clk,rst,matrix_A[12610],matrix_B[10],mul_res1[12610]);
multi_7x28 multi_7x28_mod_12611(clk,rst,matrix_A[12611],matrix_B[11],mul_res1[12611]);
multi_7x28 multi_7x28_mod_12612(clk,rst,matrix_A[12612],matrix_B[12],mul_res1[12612]);
multi_7x28 multi_7x28_mod_12613(clk,rst,matrix_A[12613],matrix_B[13],mul_res1[12613]);
multi_7x28 multi_7x28_mod_12614(clk,rst,matrix_A[12614],matrix_B[14],mul_res1[12614]);
multi_7x28 multi_7x28_mod_12615(clk,rst,matrix_A[12615],matrix_B[15],mul_res1[12615]);
multi_7x28 multi_7x28_mod_12616(clk,rst,matrix_A[12616],matrix_B[16],mul_res1[12616]);
multi_7x28 multi_7x28_mod_12617(clk,rst,matrix_A[12617],matrix_B[17],mul_res1[12617]);
multi_7x28 multi_7x28_mod_12618(clk,rst,matrix_A[12618],matrix_B[18],mul_res1[12618]);
multi_7x28 multi_7x28_mod_12619(clk,rst,matrix_A[12619],matrix_B[19],mul_res1[12619]);
multi_7x28 multi_7x28_mod_12620(clk,rst,matrix_A[12620],matrix_B[20],mul_res1[12620]);
multi_7x28 multi_7x28_mod_12621(clk,rst,matrix_A[12621],matrix_B[21],mul_res1[12621]);
multi_7x28 multi_7x28_mod_12622(clk,rst,matrix_A[12622],matrix_B[22],mul_res1[12622]);
multi_7x28 multi_7x28_mod_12623(clk,rst,matrix_A[12623],matrix_B[23],mul_res1[12623]);
multi_7x28 multi_7x28_mod_12624(clk,rst,matrix_A[12624],matrix_B[24],mul_res1[12624]);
multi_7x28 multi_7x28_mod_12625(clk,rst,matrix_A[12625],matrix_B[25],mul_res1[12625]);
multi_7x28 multi_7x28_mod_12626(clk,rst,matrix_A[12626],matrix_B[26],mul_res1[12626]);
multi_7x28 multi_7x28_mod_12627(clk,rst,matrix_A[12627],matrix_B[27],mul_res1[12627]);
multi_7x28 multi_7x28_mod_12628(clk,rst,matrix_A[12628],matrix_B[28],mul_res1[12628]);
multi_7x28 multi_7x28_mod_12629(clk,rst,matrix_A[12629],matrix_B[29],mul_res1[12629]);
multi_7x28 multi_7x28_mod_12630(clk,rst,matrix_A[12630],matrix_B[30],mul_res1[12630]);
multi_7x28 multi_7x28_mod_12631(clk,rst,matrix_A[12631],matrix_B[31],mul_res1[12631]);
multi_7x28 multi_7x28_mod_12632(clk,rst,matrix_A[12632],matrix_B[32],mul_res1[12632]);
multi_7x28 multi_7x28_mod_12633(clk,rst,matrix_A[12633],matrix_B[33],mul_res1[12633]);
multi_7x28 multi_7x28_mod_12634(clk,rst,matrix_A[12634],matrix_B[34],mul_res1[12634]);
multi_7x28 multi_7x28_mod_12635(clk,rst,matrix_A[12635],matrix_B[35],mul_res1[12635]);
multi_7x28 multi_7x28_mod_12636(clk,rst,matrix_A[12636],matrix_B[36],mul_res1[12636]);
multi_7x28 multi_7x28_mod_12637(clk,rst,matrix_A[12637],matrix_B[37],mul_res1[12637]);
multi_7x28 multi_7x28_mod_12638(clk,rst,matrix_A[12638],matrix_B[38],mul_res1[12638]);
multi_7x28 multi_7x28_mod_12639(clk,rst,matrix_A[12639],matrix_B[39],mul_res1[12639]);
multi_7x28 multi_7x28_mod_12640(clk,rst,matrix_A[12640],matrix_B[40],mul_res1[12640]);
multi_7x28 multi_7x28_mod_12641(clk,rst,matrix_A[12641],matrix_B[41],mul_res1[12641]);
multi_7x28 multi_7x28_mod_12642(clk,rst,matrix_A[12642],matrix_B[42],mul_res1[12642]);
multi_7x28 multi_7x28_mod_12643(clk,rst,matrix_A[12643],matrix_B[43],mul_res1[12643]);
multi_7x28 multi_7x28_mod_12644(clk,rst,matrix_A[12644],matrix_B[44],mul_res1[12644]);
multi_7x28 multi_7x28_mod_12645(clk,rst,matrix_A[12645],matrix_B[45],mul_res1[12645]);
multi_7x28 multi_7x28_mod_12646(clk,rst,matrix_A[12646],matrix_B[46],mul_res1[12646]);
multi_7x28 multi_7x28_mod_12647(clk,rst,matrix_A[12647],matrix_B[47],mul_res1[12647]);
multi_7x28 multi_7x28_mod_12648(clk,rst,matrix_A[12648],matrix_B[48],mul_res1[12648]);
multi_7x28 multi_7x28_mod_12649(clk,rst,matrix_A[12649],matrix_B[49],mul_res1[12649]);
multi_7x28 multi_7x28_mod_12650(clk,rst,matrix_A[12650],matrix_B[50],mul_res1[12650]);
multi_7x28 multi_7x28_mod_12651(clk,rst,matrix_A[12651],matrix_B[51],mul_res1[12651]);
multi_7x28 multi_7x28_mod_12652(clk,rst,matrix_A[12652],matrix_B[52],mul_res1[12652]);
multi_7x28 multi_7x28_mod_12653(clk,rst,matrix_A[12653],matrix_B[53],mul_res1[12653]);
multi_7x28 multi_7x28_mod_12654(clk,rst,matrix_A[12654],matrix_B[54],mul_res1[12654]);
multi_7x28 multi_7x28_mod_12655(clk,rst,matrix_A[12655],matrix_B[55],mul_res1[12655]);
multi_7x28 multi_7x28_mod_12656(clk,rst,matrix_A[12656],matrix_B[56],mul_res1[12656]);
multi_7x28 multi_7x28_mod_12657(clk,rst,matrix_A[12657],matrix_B[57],mul_res1[12657]);
multi_7x28 multi_7x28_mod_12658(clk,rst,matrix_A[12658],matrix_B[58],mul_res1[12658]);
multi_7x28 multi_7x28_mod_12659(clk,rst,matrix_A[12659],matrix_B[59],mul_res1[12659]);
multi_7x28 multi_7x28_mod_12660(clk,rst,matrix_A[12660],matrix_B[60],mul_res1[12660]);
multi_7x28 multi_7x28_mod_12661(clk,rst,matrix_A[12661],matrix_B[61],mul_res1[12661]);
multi_7x28 multi_7x28_mod_12662(clk,rst,matrix_A[12662],matrix_B[62],mul_res1[12662]);
multi_7x28 multi_7x28_mod_12663(clk,rst,matrix_A[12663],matrix_B[63],mul_res1[12663]);
multi_7x28 multi_7x28_mod_12664(clk,rst,matrix_A[12664],matrix_B[64],mul_res1[12664]);
multi_7x28 multi_7x28_mod_12665(clk,rst,matrix_A[12665],matrix_B[65],mul_res1[12665]);
multi_7x28 multi_7x28_mod_12666(clk,rst,matrix_A[12666],matrix_B[66],mul_res1[12666]);
multi_7x28 multi_7x28_mod_12667(clk,rst,matrix_A[12667],matrix_B[67],mul_res1[12667]);
multi_7x28 multi_7x28_mod_12668(clk,rst,matrix_A[12668],matrix_B[68],mul_res1[12668]);
multi_7x28 multi_7x28_mod_12669(clk,rst,matrix_A[12669],matrix_B[69],mul_res1[12669]);
multi_7x28 multi_7x28_mod_12670(clk,rst,matrix_A[12670],matrix_B[70],mul_res1[12670]);
multi_7x28 multi_7x28_mod_12671(clk,rst,matrix_A[12671],matrix_B[71],mul_res1[12671]);
multi_7x28 multi_7x28_mod_12672(clk,rst,matrix_A[12672],matrix_B[72],mul_res1[12672]);
multi_7x28 multi_7x28_mod_12673(clk,rst,matrix_A[12673],matrix_B[73],mul_res1[12673]);
multi_7x28 multi_7x28_mod_12674(clk,rst,matrix_A[12674],matrix_B[74],mul_res1[12674]);
multi_7x28 multi_7x28_mod_12675(clk,rst,matrix_A[12675],matrix_B[75],mul_res1[12675]);
multi_7x28 multi_7x28_mod_12676(clk,rst,matrix_A[12676],matrix_B[76],mul_res1[12676]);
multi_7x28 multi_7x28_mod_12677(clk,rst,matrix_A[12677],matrix_B[77],mul_res1[12677]);
multi_7x28 multi_7x28_mod_12678(clk,rst,matrix_A[12678],matrix_B[78],mul_res1[12678]);
multi_7x28 multi_7x28_mod_12679(clk,rst,matrix_A[12679],matrix_B[79],mul_res1[12679]);
multi_7x28 multi_7x28_mod_12680(clk,rst,matrix_A[12680],matrix_B[80],mul_res1[12680]);
multi_7x28 multi_7x28_mod_12681(clk,rst,matrix_A[12681],matrix_B[81],mul_res1[12681]);
multi_7x28 multi_7x28_mod_12682(clk,rst,matrix_A[12682],matrix_B[82],mul_res1[12682]);
multi_7x28 multi_7x28_mod_12683(clk,rst,matrix_A[12683],matrix_B[83],mul_res1[12683]);
multi_7x28 multi_7x28_mod_12684(clk,rst,matrix_A[12684],matrix_B[84],mul_res1[12684]);
multi_7x28 multi_7x28_mod_12685(clk,rst,matrix_A[12685],matrix_B[85],mul_res1[12685]);
multi_7x28 multi_7x28_mod_12686(clk,rst,matrix_A[12686],matrix_B[86],mul_res1[12686]);
multi_7x28 multi_7x28_mod_12687(clk,rst,matrix_A[12687],matrix_B[87],mul_res1[12687]);
multi_7x28 multi_7x28_mod_12688(clk,rst,matrix_A[12688],matrix_B[88],mul_res1[12688]);
multi_7x28 multi_7x28_mod_12689(clk,rst,matrix_A[12689],matrix_B[89],mul_res1[12689]);
multi_7x28 multi_7x28_mod_12690(clk,rst,matrix_A[12690],matrix_B[90],mul_res1[12690]);
multi_7x28 multi_7x28_mod_12691(clk,rst,matrix_A[12691],matrix_B[91],mul_res1[12691]);
multi_7x28 multi_7x28_mod_12692(clk,rst,matrix_A[12692],matrix_B[92],mul_res1[12692]);
multi_7x28 multi_7x28_mod_12693(clk,rst,matrix_A[12693],matrix_B[93],mul_res1[12693]);
multi_7x28 multi_7x28_mod_12694(clk,rst,matrix_A[12694],matrix_B[94],mul_res1[12694]);
multi_7x28 multi_7x28_mod_12695(clk,rst,matrix_A[12695],matrix_B[95],mul_res1[12695]);
multi_7x28 multi_7x28_mod_12696(clk,rst,matrix_A[12696],matrix_B[96],mul_res1[12696]);
multi_7x28 multi_7x28_mod_12697(clk,rst,matrix_A[12697],matrix_B[97],mul_res1[12697]);
multi_7x28 multi_7x28_mod_12698(clk,rst,matrix_A[12698],matrix_B[98],mul_res1[12698]);
multi_7x28 multi_7x28_mod_12699(clk,rst,matrix_A[12699],matrix_B[99],mul_res1[12699]);
multi_7x28 multi_7x28_mod_12700(clk,rst,matrix_A[12700],matrix_B[100],mul_res1[12700]);
multi_7x28 multi_7x28_mod_12701(clk,rst,matrix_A[12701],matrix_B[101],mul_res1[12701]);
multi_7x28 multi_7x28_mod_12702(clk,rst,matrix_A[12702],matrix_B[102],mul_res1[12702]);
multi_7x28 multi_7x28_mod_12703(clk,rst,matrix_A[12703],matrix_B[103],mul_res1[12703]);
multi_7x28 multi_7x28_mod_12704(clk,rst,matrix_A[12704],matrix_B[104],mul_res1[12704]);
multi_7x28 multi_7x28_mod_12705(clk,rst,matrix_A[12705],matrix_B[105],mul_res1[12705]);
multi_7x28 multi_7x28_mod_12706(clk,rst,matrix_A[12706],matrix_B[106],mul_res1[12706]);
multi_7x28 multi_7x28_mod_12707(clk,rst,matrix_A[12707],matrix_B[107],mul_res1[12707]);
multi_7x28 multi_7x28_mod_12708(clk,rst,matrix_A[12708],matrix_B[108],mul_res1[12708]);
multi_7x28 multi_7x28_mod_12709(clk,rst,matrix_A[12709],matrix_B[109],mul_res1[12709]);
multi_7x28 multi_7x28_mod_12710(clk,rst,matrix_A[12710],matrix_B[110],mul_res1[12710]);
multi_7x28 multi_7x28_mod_12711(clk,rst,matrix_A[12711],matrix_B[111],mul_res1[12711]);
multi_7x28 multi_7x28_mod_12712(clk,rst,matrix_A[12712],matrix_B[112],mul_res1[12712]);
multi_7x28 multi_7x28_mod_12713(clk,rst,matrix_A[12713],matrix_B[113],mul_res1[12713]);
multi_7x28 multi_7x28_mod_12714(clk,rst,matrix_A[12714],matrix_B[114],mul_res1[12714]);
multi_7x28 multi_7x28_mod_12715(clk,rst,matrix_A[12715],matrix_B[115],mul_res1[12715]);
multi_7x28 multi_7x28_mod_12716(clk,rst,matrix_A[12716],matrix_B[116],mul_res1[12716]);
multi_7x28 multi_7x28_mod_12717(clk,rst,matrix_A[12717],matrix_B[117],mul_res1[12717]);
multi_7x28 multi_7x28_mod_12718(clk,rst,matrix_A[12718],matrix_B[118],mul_res1[12718]);
multi_7x28 multi_7x28_mod_12719(clk,rst,matrix_A[12719],matrix_B[119],mul_res1[12719]);
multi_7x28 multi_7x28_mod_12720(clk,rst,matrix_A[12720],matrix_B[120],mul_res1[12720]);
multi_7x28 multi_7x28_mod_12721(clk,rst,matrix_A[12721],matrix_B[121],mul_res1[12721]);
multi_7x28 multi_7x28_mod_12722(clk,rst,matrix_A[12722],matrix_B[122],mul_res1[12722]);
multi_7x28 multi_7x28_mod_12723(clk,rst,matrix_A[12723],matrix_B[123],mul_res1[12723]);
multi_7x28 multi_7x28_mod_12724(clk,rst,matrix_A[12724],matrix_B[124],mul_res1[12724]);
multi_7x28 multi_7x28_mod_12725(clk,rst,matrix_A[12725],matrix_B[125],mul_res1[12725]);
multi_7x28 multi_7x28_mod_12726(clk,rst,matrix_A[12726],matrix_B[126],mul_res1[12726]);
multi_7x28 multi_7x28_mod_12727(clk,rst,matrix_A[12727],matrix_B[127],mul_res1[12727]);
multi_7x28 multi_7x28_mod_12728(clk,rst,matrix_A[12728],matrix_B[128],mul_res1[12728]);
multi_7x28 multi_7x28_mod_12729(clk,rst,matrix_A[12729],matrix_B[129],mul_res1[12729]);
multi_7x28 multi_7x28_mod_12730(clk,rst,matrix_A[12730],matrix_B[130],mul_res1[12730]);
multi_7x28 multi_7x28_mod_12731(clk,rst,matrix_A[12731],matrix_B[131],mul_res1[12731]);
multi_7x28 multi_7x28_mod_12732(clk,rst,matrix_A[12732],matrix_B[132],mul_res1[12732]);
multi_7x28 multi_7x28_mod_12733(clk,rst,matrix_A[12733],matrix_B[133],mul_res1[12733]);
multi_7x28 multi_7x28_mod_12734(clk,rst,matrix_A[12734],matrix_B[134],mul_res1[12734]);
multi_7x28 multi_7x28_mod_12735(clk,rst,matrix_A[12735],matrix_B[135],mul_res1[12735]);
multi_7x28 multi_7x28_mod_12736(clk,rst,matrix_A[12736],matrix_B[136],mul_res1[12736]);
multi_7x28 multi_7x28_mod_12737(clk,rst,matrix_A[12737],matrix_B[137],mul_res1[12737]);
multi_7x28 multi_7x28_mod_12738(clk,rst,matrix_A[12738],matrix_B[138],mul_res1[12738]);
multi_7x28 multi_7x28_mod_12739(clk,rst,matrix_A[12739],matrix_B[139],mul_res1[12739]);
multi_7x28 multi_7x28_mod_12740(clk,rst,matrix_A[12740],matrix_B[140],mul_res1[12740]);
multi_7x28 multi_7x28_mod_12741(clk,rst,matrix_A[12741],matrix_B[141],mul_res1[12741]);
multi_7x28 multi_7x28_mod_12742(clk,rst,matrix_A[12742],matrix_B[142],mul_res1[12742]);
multi_7x28 multi_7x28_mod_12743(clk,rst,matrix_A[12743],matrix_B[143],mul_res1[12743]);
multi_7x28 multi_7x28_mod_12744(clk,rst,matrix_A[12744],matrix_B[144],mul_res1[12744]);
multi_7x28 multi_7x28_mod_12745(clk,rst,matrix_A[12745],matrix_B[145],mul_res1[12745]);
multi_7x28 multi_7x28_mod_12746(clk,rst,matrix_A[12746],matrix_B[146],mul_res1[12746]);
multi_7x28 multi_7x28_mod_12747(clk,rst,matrix_A[12747],matrix_B[147],mul_res1[12747]);
multi_7x28 multi_7x28_mod_12748(clk,rst,matrix_A[12748],matrix_B[148],mul_res1[12748]);
multi_7x28 multi_7x28_mod_12749(clk,rst,matrix_A[12749],matrix_B[149],mul_res1[12749]);
multi_7x28 multi_7x28_mod_12750(clk,rst,matrix_A[12750],matrix_B[150],mul_res1[12750]);
multi_7x28 multi_7x28_mod_12751(clk,rst,matrix_A[12751],matrix_B[151],mul_res1[12751]);
multi_7x28 multi_7x28_mod_12752(clk,rst,matrix_A[12752],matrix_B[152],mul_res1[12752]);
multi_7x28 multi_7x28_mod_12753(clk,rst,matrix_A[12753],matrix_B[153],mul_res1[12753]);
multi_7x28 multi_7x28_mod_12754(clk,rst,matrix_A[12754],matrix_B[154],mul_res1[12754]);
multi_7x28 multi_7x28_mod_12755(clk,rst,matrix_A[12755],matrix_B[155],mul_res1[12755]);
multi_7x28 multi_7x28_mod_12756(clk,rst,matrix_A[12756],matrix_B[156],mul_res1[12756]);
multi_7x28 multi_7x28_mod_12757(clk,rst,matrix_A[12757],matrix_B[157],mul_res1[12757]);
multi_7x28 multi_7x28_mod_12758(clk,rst,matrix_A[12758],matrix_B[158],mul_res1[12758]);
multi_7x28 multi_7x28_mod_12759(clk,rst,matrix_A[12759],matrix_B[159],mul_res1[12759]);
multi_7x28 multi_7x28_mod_12760(clk,rst,matrix_A[12760],matrix_B[160],mul_res1[12760]);
multi_7x28 multi_7x28_mod_12761(clk,rst,matrix_A[12761],matrix_B[161],mul_res1[12761]);
multi_7x28 multi_7x28_mod_12762(clk,rst,matrix_A[12762],matrix_B[162],mul_res1[12762]);
multi_7x28 multi_7x28_mod_12763(clk,rst,matrix_A[12763],matrix_B[163],mul_res1[12763]);
multi_7x28 multi_7x28_mod_12764(clk,rst,matrix_A[12764],matrix_B[164],mul_res1[12764]);
multi_7x28 multi_7x28_mod_12765(clk,rst,matrix_A[12765],matrix_B[165],mul_res1[12765]);
multi_7x28 multi_7x28_mod_12766(clk,rst,matrix_A[12766],matrix_B[166],mul_res1[12766]);
multi_7x28 multi_7x28_mod_12767(clk,rst,matrix_A[12767],matrix_B[167],mul_res1[12767]);
multi_7x28 multi_7x28_mod_12768(clk,rst,matrix_A[12768],matrix_B[168],mul_res1[12768]);
multi_7x28 multi_7x28_mod_12769(clk,rst,matrix_A[12769],matrix_B[169],mul_res1[12769]);
multi_7x28 multi_7x28_mod_12770(clk,rst,matrix_A[12770],matrix_B[170],mul_res1[12770]);
multi_7x28 multi_7x28_mod_12771(clk,rst,matrix_A[12771],matrix_B[171],mul_res1[12771]);
multi_7x28 multi_7x28_mod_12772(clk,rst,matrix_A[12772],matrix_B[172],mul_res1[12772]);
multi_7x28 multi_7x28_mod_12773(clk,rst,matrix_A[12773],matrix_B[173],mul_res1[12773]);
multi_7x28 multi_7x28_mod_12774(clk,rst,matrix_A[12774],matrix_B[174],mul_res1[12774]);
multi_7x28 multi_7x28_mod_12775(clk,rst,matrix_A[12775],matrix_B[175],mul_res1[12775]);
multi_7x28 multi_7x28_mod_12776(clk,rst,matrix_A[12776],matrix_B[176],mul_res1[12776]);
multi_7x28 multi_7x28_mod_12777(clk,rst,matrix_A[12777],matrix_B[177],mul_res1[12777]);
multi_7x28 multi_7x28_mod_12778(clk,rst,matrix_A[12778],matrix_B[178],mul_res1[12778]);
multi_7x28 multi_7x28_mod_12779(clk,rst,matrix_A[12779],matrix_B[179],mul_res1[12779]);
multi_7x28 multi_7x28_mod_12780(clk,rst,matrix_A[12780],matrix_B[180],mul_res1[12780]);
multi_7x28 multi_7x28_mod_12781(clk,rst,matrix_A[12781],matrix_B[181],mul_res1[12781]);
multi_7x28 multi_7x28_mod_12782(clk,rst,matrix_A[12782],matrix_B[182],mul_res1[12782]);
multi_7x28 multi_7x28_mod_12783(clk,rst,matrix_A[12783],matrix_B[183],mul_res1[12783]);
multi_7x28 multi_7x28_mod_12784(clk,rst,matrix_A[12784],matrix_B[184],mul_res1[12784]);
multi_7x28 multi_7x28_mod_12785(clk,rst,matrix_A[12785],matrix_B[185],mul_res1[12785]);
multi_7x28 multi_7x28_mod_12786(clk,rst,matrix_A[12786],matrix_B[186],mul_res1[12786]);
multi_7x28 multi_7x28_mod_12787(clk,rst,matrix_A[12787],matrix_B[187],mul_res1[12787]);
multi_7x28 multi_7x28_mod_12788(clk,rst,matrix_A[12788],matrix_B[188],mul_res1[12788]);
multi_7x28 multi_7x28_mod_12789(clk,rst,matrix_A[12789],matrix_B[189],mul_res1[12789]);
multi_7x28 multi_7x28_mod_12790(clk,rst,matrix_A[12790],matrix_B[190],mul_res1[12790]);
multi_7x28 multi_7x28_mod_12791(clk,rst,matrix_A[12791],matrix_B[191],mul_res1[12791]);
multi_7x28 multi_7x28_mod_12792(clk,rst,matrix_A[12792],matrix_B[192],mul_res1[12792]);
multi_7x28 multi_7x28_mod_12793(clk,rst,matrix_A[12793],matrix_B[193],mul_res1[12793]);
multi_7x28 multi_7x28_mod_12794(clk,rst,matrix_A[12794],matrix_B[194],mul_res1[12794]);
multi_7x28 multi_7x28_mod_12795(clk,rst,matrix_A[12795],matrix_B[195],mul_res1[12795]);
multi_7x28 multi_7x28_mod_12796(clk,rst,matrix_A[12796],matrix_B[196],mul_res1[12796]);
multi_7x28 multi_7x28_mod_12797(clk,rst,matrix_A[12797],matrix_B[197],mul_res1[12797]);
multi_7x28 multi_7x28_mod_12798(clk,rst,matrix_A[12798],matrix_B[198],mul_res1[12798]);
multi_7x28 multi_7x28_mod_12799(clk,rst,matrix_A[12799],matrix_B[199],mul_res1[12799]);
 
 
 
 
/*


#include <stdio.h>
   
   int main() {
       // Write C code here
       int i,j;
       int k = 0;
       int z = 0;
      for (i = 0; i<=63; i++) { //64-1
        for (j = 0; j<= 199;j++) {     //200-1
          z = ((64 * j) - 1 + i) < 0 ? 0 : ((64 * j)  + i); // 64 is width of matrix
printf("multi_7x28 multi_7x28_mod_%d(clk,rst,matrix_A[%d],matrix_B[%d],mul_res1[%d]);\n",k,k,j,k);
k = k+1;
}
}
       return 0;
   }

*/

adder_200in adder_200in_mod_0(clk,rst,mul_res1[0],mul_res1[1],mul_res1[2],mul_res1[3],mul_res1[4],mul_res1[5],mul_res1[6],mul_res1[7],mul_res1[8],mul_res1[9],mul_res1[10],mul_res1[11],mul_res1[12],mul_res1[13],mul_res1[14],mul_res1[15],mul_res1[16],mul_res1[17],mul_res1[18],mul_res1[19],mul_res1[20],mul_res1[21],mul_res1[22],mul_res1[23],mul_res1[24],mul_res1[25],mul_res1[26],mul_res1[27],mul_res1[28],mul_res1[29],mul_res1[30],mul_res1[31],mul_res1[32],mul_res1[33],mul_res1[34],mul_res1[35],mul_res1[36],mul_res1[37],mul_res1[38],mul_res1[39],mul_res1[40],mul_res1[41],mul_res1[42],mul_res1[43],mul_res1[44],mul_res1[45],mul_res1[46],mul_res1[47],mul_res1[48],mul_res1[49],mul_res1[50],mul_res1[51],mul_res1[52],mul_res1[53],mul_res1[54],mul_res1[55],mul_res1[56],mul_res1[57],mul_res1[58],mul_res1[59],mul_res1[60],mul_res1[61],mul_res1[62],mul_res1[63],mul_res1[64],mul_res1[65],mul_res1[66],mul_res1[67],mul_res1[68],mul_res1[69],mul_res1[70],mul_res1[71],mul_res1[72],mul_res1[73],mul_res1[74],mul_res1[75],mul_res1[76],mul_res1[77],mul_res1[78],mul_res1[79],mul_res1[80],mul_res1[81],mul_res1[82],mul_res1[83],mul_res1[84],mul_res1[85],mul_res1[86],mul_res1[87],mul_res1[88],mul_res1[89],mul_res1[90],mul_res1[91],mul_res1[92],mul_res1[93],mul_res1[94],mul_res1[95],mul_res1[96],mul_res1[97],mul_res1[98],mul_res1[99],mul_res1[100],mul_res1[101],mul_res1[102],mul_res1[103],mul_res1[104],mul_res1[105],mul_res1[106],mul_res1[107],mul_res1[108],mul_res1[109],mul_res1[110],mul_res1[111],mul_res1[112],mul_res1[113],mul_res1[114],mul_res1[115],mul_res1[116],mul_res1[117],mul_res1[118],mul_res1[119],mul_res1[120],mul_res1[121],mul_res1[122],mul_res1[123],mul_res1[124],mul_res1[125],mul_res1[126],mul_res1[127],mul_res1[128],mul_res1[129],mul_res1[130],mul_res1[131],mul_res1[132],mul_res1[133],mul_res1[134],mul_res1[135],mul_res1[136],mul_res1[137],mul_res1[138],mul_res1[139],mul_res1[140],mul_res1[141],mul_res1[142],mul_res1[143],mul_res1[144],mul_res1[145],mul_res1[146],mul_res1[147],mul_res1[148],mul_res1[149],mul_res1[150],mul_res1[151],mul_res1[152],mul_res1[153],mul_res1[154],mul_res1[155],mul_res1[156],mul_res1[157],mul_res1[158],mul_res1[159],mul_res1[160],mul_res1[161],mul_res1[162],mul_res1[163],mul_res1[164],mul_res1[165],mul_res1[166],mul_res1[167],mul_res1[168],mul_res1[169],mul_res1[170],mul_res1[171],mul_res1[172],mul_res1[173],mul_res1[174],mul_res1[175],mul_res1[176],mul_res1[177],mul_res1[178],mul_res1[179],mul_res1[180],mul_res1[181],mul_res1[182],mul_res1[183],mul_res1[184],mul_res1[185],mul_res1[186],mul_res1[187],mul_res1[188],mul_res1[189],mul_res1[190],mul_res1[191],mul_res1[192],mul_res1[193],mul_res1[194],mul_res1[195],mul_res1[196],mul_res1[197],mul_res1[198],mul_res1[199],result_fc1[0]);


adder_200in adder_200in_mod_1(clk,rst,mul_res1[200],mul_res1[201],mul_res1[202],mul_res1[203],mul_res1[204],mul_res1[205],mul_res1[206],mul_res1[207],mul_res1[208],mul_res1[209],mul_res1[210],mul_res1[211],mul_res1[212],mul_res1[213],mul_res1[214],mul_res1[215],mul_res1[216],mul_res1[217],mul_res1[218],mul_res1[219],mul_res1[220],mul_res1[221],mul_res1[222],mul_res1[223],mul_res1[224],mul_res1[225],mul_res1[226],mul_res1[227],mul_res1[228],mul_res1[229],mul_res1[230],mul_res1[231],mul_res1[232],mul_res1[233],mul_res1[234],mul_res1[235],mul_res1[236],mul_res1[237],mul_res1[238],mul_res1[239],mul_res1[240],mul_res1[241],mul_res1[242],mul_res1[243],mul_res1[244],mul_res1[245],mul_res1[246],mul_res1[247],mul_res1[248],mul_res1[249],mul_res1[250],mul_res1[251],mul_res1[252],mul_res1[253],mul_res1[254],mul_res1[255],mul_res1[256],mul_res1[257],mul_res1[258],mul_res1[259],mul_res1[260],mul_res1[261],mul_res1[262],mul_res1[263],mul_res1[264],mul_res1[265],mul_res1[266],mul_res1[267],mul_res1[268],mul_res1[269],mul_res1[270],mul_res1[271],mul_res1[272],mul_res1[273],mul_res1[274],mul_res1[275],mul_res1[276],mul_res1[277],mul_res1[278],mul_res1[279],mul_res1[280],mul_res1[281],mul_res1[282],mul_res1[283],mul_res1[284],mul_res1[285],mul_res1[286],mul_res1[287],mul_res1[288],mul_res1[289],mul_res1[290],mul_res1[291],mul_res1[292],mul_res1[293],mul_res1[294],mul_res1[295],mul_res1[296],mul_res1[297],mul_res1[298],mul_res1[299],mul_res1[300],mul_res1[301],mul_res1[302],mul_res1[303],mul_res1[304],mul_res1[305],mul_res1[306],mul_res1[307],mul_res1[308],mul_res1[309],mul_res1[310],mul_res1[311],mul_res1[312],mul_res1[313],mul_res1[314],mul_res1[315],mul_res1[316],mul_res1[317],mul_res1[318],mul_res1[319],mul_res1[320],mul_res1[321],mul_res1[322],mul_res1[323],mul_res1[324],mul_res1[325],mul_res1[326],mul_res1[327],mul_res1[328],mul_res1[329],mul_res1[330],mul_res1[331],mul_res1[332],mul_res1[333],mul_res1[334],mul_res1[335],mul_res1[336],mul_res1[337],mul_res1[338],mul_res1[339],mul_res1[340],mul_res1[341],mul_res1[342],mul_res1[343],mul_res1[344],mul_res1[345],mul_res1[346],mul_res1[347],mul_res1[348],mul_res1[349],mul_res1[350],mul_res1[351],mul_res1[352],mul_res1[353],mul_res1[354],mul_res1[355],mul_res1[356],mul_res1[357],mul_res1[358],mul_res1[359],mul_res1[360],mul_res1[361],mul_res1[362],mul_res1[363],mul_res1[364],mul_res1[365],mul_res1[366],mul_res1[367],mul_res1[368],mul_res1[369],mul_res1[370],mul_res1[371],mul_res1[372],mul_res1[373],mul_res1[374],mul_res1[375],mul_res1[376],mul_res1[377],mul_res1[378],mul_res1[379],mul_res1[380],mul_res1[381],mul_res1[382],mul_res1[383],mul_res1[384],mul_res1[385],mul_res1[386],mul_res1[387],mul_res1[388],mul_res1[389],mul_res1[390],mul_res1[391],mul_res1[392],mul_res1[393],mul_res1[394],mul_res1[395],mul_res1[396],mul_res1[397],mul_res1[398],mul_res1[399],result_fc1[1]);


adder_200in adder_200in_mod_2(clk,rst,mul_res1[400],mul_res1[401],mul_res1[402],mul_res1[403],mul_res1[404],mul_res1[405],mul_res1[406],mul_res1[407],mul_res1[408],mul_res1[409],mul_res1[410],mul_res1[411],mul_res1[412],mul_res1[413],mul_res1[414],mul_res1[415],mul_res1[416],mul_res1[417],mul_res1[418],mul_res1[419],mul_res1[420],mul_res1[421],mul_res1[422],mul_res1[423],mul_res1[424],mul_res1[425],mul_res1[426],mul_res1[427],mul_res1[428],mul_res1[429],mul_res1[430],mul_res1[431],mul_res1[432],mul_res1[433],mul_res1[434],mul_res1[435],mul_res1[436],mul_res1[437],mul_res1[438],mul_res1[439],mul_res1[440],mul_res1[441],mul_res1[442],mul_res1[443],mul_res1[444],mul_res1[445],mul_res1[446],mul_res1[447],mul_res1[448],mul_res1[449],mul_res1[450],mul_res1[451],mul_res1[452],mul_res1[453],mul_res1[454],mul_res1[455],mul_res1[456],mul_res1[457],mul_res1[458],mul_res1[459],mul_res1[460],mul_res1[461],mul_res1[462],mul_res1[463],mul_res1[464],mul_res1[465],mul_res1[466],mul_res1[467],mul_res1[468],mul_res1[469],mul_res1[470],mul_res1[471],mul_res1[472],mul_res1[473],mul_res1[474],mul_res1[475],mul_res1[476],mul_res1[477],mul_res1[478],mul_res1[479],mul_res1[480],mul_res1[481],mul_res1[482],mul_res1[483],mul_res1[484],mul_res1[485],mul_res1[486],mul_res1[487],mul_res1[488],mul_res1[489],mul_res1[490],mul_res1[491],mul_res1[492],mul_res1[493],mul_res1[494],mul_res1[495],mul_res1[496],mul_res1[497],mul_res1[498],mul_res1[499],mul_res1[500],mul_res1[501],mul_res1[502],mul_res1[503],mul_res1[504],mul_res1[505],mul_res1[506],mul_res1[507],mul_res1[508],mul_res1[509],mul_res1[510],mul_res1[511],mul_res1[512],mul_res1[513],mul_res1[514],mul_res1[515],mul_res1[516],mul_res1[517],mul_res1[518],mul_res1[519],mul_res1[520],mul_res1[521],mul_res1[522],mul_res1[523],mul_res1[524],mul_res1[525],mul_res1[526],mul_res1[527],mul_res1[528],mul_res1[529],mul_res1[530],mul_res1[531],mul_res1[532],mul_res1[533],mul_res1[534],mul_res1[535],mul_res1[536],mul_res1[537],mul_res1[538],mul_res1[539],mul_res1[540],mul_res1[541],mul_res1[542],mul_res1[543],mul_res1[544],mul_res1[545],mul_res1[546],mul_res1[547],mul_res1[548],mul_res1[549],mul_res1[550],mul_res1[551],mul_res1[552],mul_res1[553],mul_res1[554],mul_res1[555],mul_res1[556],mul_res1[557],mul_res1[558],mul_res1[559],mul_res1[560],mul_res1[561],mul_res1[562],mul_res1[563],mul_res1[564],mul_res1[565],mul_res1[566],mul_res1[567],mul_res1[568],mul_res1[569],mul_res1[570],mul_res1[571],mul_res1[572],mul_res1[573],mul_res1[574],mul_res1[575],mul_res1[576],mul_res1[577],mul_res1[578],mul_res1[579],mul_res1[580],mul_res1[581],mul_res1[582],mul_res1[583],mul_res1[584],mul_res1[585],mul_res1[586],mul_res1[587],mul_res1[588],mul_res1[589],mul_res1[590],mul_res1[591],mul_res1[592],mul_res1[593],mul_res1[594],mul_res1[595],mul_res1[596],mul_res1[597],mul_res1[598],mul_res1[599],result_fc1[2]);


adder_200in adder_200in_mod_3(clk,rst,mul_res1[600],mul_res1[601],mul_res1[602],mul_res1[603],mul_res1[604],mul_res1[605],mul_res1[606],mul_res1[607],mul_res1[608],mul_res1[609],mul_res1[610],mul_res1[611],mul_res1[612],mul_res1[613],mul_res1[614],mul_res1[615],mul_res1[616],mul_res1[617],mul_res1[618],mul_res1[619],mul_res1[620],mul_res1[621],mul_res1[622],mul_res1[623],mul_res1[624],mul_res1[625],mul_res1[626],mul_res1[627],mul_res1[628],mul_res1[629],mul_res1[630],mul_res1[631],mul_res1[632],mul_res1[633],mul_res1[634],mul_res1[635],mul_res1[636],mul_res1[637],mul_res1[638],mul_res1[639],mul_res1[640],mul_res1[641],mul_res1[642],mul_res1[643],mul_res1[644],mul_res1[645],mul_res1[646],mul_res1[647],mul_res1[648],mul_res1[649],mul_res1[650],mul_res1[651],mul_res1[652],mul_res1[653],mul_res1[654],mul_res1[655],mul_res1[656],mul_res1[657],mul_res1[658],mul_res1[659],mul_res1[660],mul_res1[661],mul_res1[662],mul_res1[663],mul_res1[664],mul_res1[665],mul_res1[666],mul_res1[667],mul_res1[668],mul_res1[669],mul_res1[670],mul_res1[671],mul_res1[672],mul_res1[673],mul_res1[674],mul_res1[675],mul_res1[676],mul_res1[677],mul_res1[678],mul_res1[679],mul_res1[680],mul_res1[681],mul_res1[682],mul_res1[683],mul_res1[684],mul_res1[685],mul_res1[686],mul_res1[687],mul_res1[688],mul_res1[689],mul_res1[690],mul_res1[691],mul_res1[692],mul_res1[693],mul_res1[694],mul_res1[695],mul_res1[696],mul_res1[697],mul_res1[698],mul_res1[699],mul_res1[700],mul_res1[701],mul_res1[702],mul_res1[703],mul_res1[704],mul_res1[705],mul_res1[706],mul_res1[707],mul_res1[708],mul_res1[709],mul_res1[710],mul_res1[711],mul_res1[712],mul_res1[713],mul_res1[714],mul_res1[715],mul_res1[716],mul_res1[717],mul_res1[718],mul_res1[719],mul_res1[720],mul_res1[721],mul_res1[722],mul_res1[723],mul_res1[724],mul_res1[725],mul_res1[726],mul_res1[727],mul_res1[728],mul_res1[729],mul_res1[730],mul_res1[731],mul_res1[732],mul_res1[733],mul_res1[734],mul_res1[735],mul_res1[736],mul_res1[737],mul_res1[738],mul_res1[739],mul_res1[740],mul_res1[741],mul_res1[742],mul_res1[743],mul_res1[744],mul_res1[745],mul_res1[746],mul_res1[747],mul_res1[748],mul_res1[749],mul_res1[750],mul_res1[751],mul_res1[752],mul_res1[753],mul_res1[754],mul_res1[755],mul_res1[756],mul_res1[757],mul_res1[758],mul_res1[759],mul_res1[760],mul_res1[761],mul_res1[762],mul_res1[763],mul_res1[764],mul_res1[765],mul_res1[766],mul_res1[767],mul_res1[768],mul_res1[769],mul_res1[770],mul_res1[771],mul_res1[772],mul_res1[773],mul_res1[774],mul_res1[775],mul_res1[776],mul_res1[777],mul_res1[778],mul_res1[779],mul_res1[780],mul_res1[781],mul_res1[782],mul_res1[783],mul_res1[784],mul_res1[785],mul_res1[786],mul_res1[787],mul_res1[788],mul_res1[789],mul_res1[790],mul_res1[791],mul_res1[792],mul_res1[793],mul_res1[794],mul_res1[795],mul_res1[796],mul_res1[797],mul_res1[798],mul_res1[799],result_fc1[3]);


adder_200in adder_200in_mod_4(clk,rst,mul_res1[800],mul_res1[801],mul_res1[802],mul_res1[803],mul_res1[804],mul_res1[805],mul_res1[806],mul_res1[807],mul_res1[808],mul_res1[809],mul_res1[810],mul_res1[811],mul_res1[812],mul_res1[813],mul_res1[814],mul_res1[815],mul_res1[816],mul_res1[817],mul_res1[818],mul_res1[819],mul_res1[820],mul_res1[821],mul_res1[822],mul_res1[823],mul_res1[824],mul_res1[825],mul_res1[826],mul_res1[827],mul_res1[828],mul_res1[829],mul_res1[830],mul_res1[831],mul_res1[832],mul_res1[833],mul_res1[834],mul_res1[835],mul_res1[836],mul_res1[837],mul_res1[838],mul_res1[839],mul_res1[840],mul_res1[841],mul_res1[842],mul_res1[843],mul_res1[844],mul_res1[845],mul_res1[846],mul_res1[847],mul_res1[848],mul_res1[849],mul_res1[850],mul_res1[851],mul_res1[852],mul_res1[853],mul_res1[854],mul_res1[855],mul_res1[856],mul_res1[857],mul_res1[858],mul_res1[859],mul_res1[860],mul_res1[861],mul_res1[862],mul_res1[863],mul_res1[864],mul_res1[865],mul_res1[866],mul_res1[867],mul_res1[868],mul_res1[869],mul_res1[870],mul_res1[871],mul_res1[872],mul_res1[873],mul_res1[874],mul_res1[875],mul_res1[876],mul_res1[877],mul_res1[878],mul_res1[879],mul_res1[880],mul_res1[881],mul_res1[882],mul_res1[883],mul_res1[884],mul_res1[885],mul_res1[886],mul_res1[887],mul_res1[888],mul_res1[889],mul_res1[890],mul_res1[891],mul_res1[892],mul_res1[893],mul_res1[894],mul_res1[895],mul_res1[896],mul_res1[897],mul_res1[898],mul_res1[899],mul_res1[900],mul_res1[901],mul_res1[902],mul_res1[903],mul_res1[904],mul_res1[905],mul_res1[906],mul_res1[907],mul_res1[908],mul_res1[909],mul_res1[910],mul_res1[911],mul_res1[912],mul_res1[913],mul_res1[914],mul_res1[915],mul_res1[916],mul_res1[917],mul_res1[918],mul_res1[919],mul_res1[920],mul_res1[921],mul_res1[922],mul_res1[923],mul_res1[924],mul_res1[925],mul_res1[926],mul_res1[927],mul_res1[928],mul_res1[929],mul_res1[930],mul_res1[931],mul_res1[932],mul_res1[933],mul_res1[934],mul_res1[935],mul_res1[936],mul_res1[937],mul_res1[938],mul_res1[939],mul_res1[940],mul_res1[941],mul_res1[942],mul_res1[943],mul_res1[944],mul_res1[945],mul_res1[946],mul_res1[947],mul_res1[948],mul_res1[949],mul_res1[950],mul_res1[951],mul_res1[952],mul_res1[953],mul_res1[954],mul_res1[955],mul_res1[956],mul_res1[957],mul_res1[958],mul_res1[959],mul_res1[960],mul_res1[961],mul_res1[962],mul_res1[963],mul_res1[964],mul_res1[965],mul_res1[966],mul_res1[967],mul_res1[968],mul_res1[969],mul_res1[970],mul_res1[971],mul_res1[972],mul_res1[973],mul_res1[974],mul_res1[975],mul_res1[976],mul_res1[977],mul_res1[978],mul_res1[979],mul_res1[980],mul_res1[981],mul_res1[982],mul_res1[983],mul_res1[984],mul_res1[985],mul_res1[986],mul_res1[987],mul_res1[988],mul_res1[989],mul_res1[990],mul_res1[991],mul_res1[992],mul_res1[993],mul_res1[994],mul_res1[995],mul_res1[996],mul_res1[997],mul_res1[998],mul_res1[999],result_fc1[4]);


adder_200in adder_200in_mod_5(clk,rst,mul_res1[1000],mul_res1[1001],mul_res1[1002],mul_res1[1003],mul_res1[1004],mul_res1[1005],mul_res1[1006],mul_res1[1007],mul_res1[1008],mul_res1[1009],mul_res1[1010],mul_res1[1011],mul_res1[1012],mul_res1[1013],mul_res1[1014],mul_res1[1015],mul_res1[1016],mul_res1[1017],mul_res1[1018],mul_res1[1019],mul_res1[1020],mul_res1[1021],mul_res1[1022],mul_res1[1023],mul_res1[1024],mul_res1[1025],mul_res1[1026],mul_res1[1027],mul_res1[1028],mul_res1[1029],mul_res1[1030],mul_res1[1031],mul_res1[1032],mul_res1[1033],mul_res1[1034],mul_res1[1035],mul_res1[1036],mul_res1[1037],mul_res1[1038],mul_res1[1039],mul_res1[1040],mul_res1[1041],mul_res1[1042],mul_res1[1043],mul_res1[1044],mul_res1[1045],mul_res1[1046],mul_res1[1047],mul_res1[1048],mul_res1[1049],mul_res1[1050],mul_res1[1051],mul_res1[1052],mul_res1[1053],mul_res1[1054],mul_res1[1055],mul_res1[1056],mul_res1[1057],mul_res1[1058],mul_res1[1059],mul_res1[1060],mul_res1[1061],mul_res1[1062],mul_res1[1063],mul_res1[1064],mul_res1[1065],mul_res1[1066],mul_res1[1067],mul_res1[1068],mul_res1[1069],mul_res1[1070],mul_res1[1071],mul_res1[1072],mul_res1[1073],mul_res1[1074],mul_res1[1075],mul_res1[1076],mul_res1[1077],mul_res1[1078],mul_res1[1079],mul_res1[1080],mul_res1[1081],mul_res1[1082],mul_res1[1083],mul_res1[1084],mul_res1[1085],mul_res1[1086],mul_res1[1087],mul_res1[1088],mul_res1[1089],mul_res1[1090],mul_res1[1091],mul_res1[1092],mul_res1[1093],mul_res1[1094],mul_res1[1095],mul_res1[1096],mul_res1[1097],mul_res1[1098],mul_res1[1099],mul_res1[1100],mul_res1[1101],mul_res1[1102],mul_res1[1103],mul_res1[1104],mul_res1[1105],mul_res1[1106],mul_res1[1107],mul_res1[1108],mul_res1[1109],mul_res1[1110],mul_res1[1111],mul_res1[1112],mul_res1[1113],mul_res1[1114],mul_res1[1115],mul_res1[1116],mul_res1[1117],mul_res1[1118],mul_res1[1119],mul_res1[1120],mul_res1[1121],mul_res1[1122],mul_res1[1123],mul_res1[1124],mul_res1[1125],mul_res1[1126],mul_res1[1127],mul_res1[1128],mul_res1[1129],mul_res1[1130],mul_res1[1131],mul_res1[1132],mul_res1[1133],mul_res1[1134],mul_res1[1135],mul_res1[1136],mul_res1[1137],mul_res1[1138],mul_res1[1139],mul_res1[1140],mul_res1[1141],mul_res1[1142],mul_res1[1143],mul_res1[1144],mul_res1[1145],mul_res1[1146],mul_res1[1147],mul_res1[1148],mul_res1[1149],mul_res1[1150],mul_res1[1151],mul_res1[1152],mul_res1[1153],mul_res1[1154],mul_res1[1155],mul_res1[1156],mul_res1[1157],mul_res1[1158],mul_res1[1159],mul_res1[1160],mul_res1[1161],mul_res1[1162],mul_res1[1163],mul_res1[1164],mul_res1[1165],mul_res1[1166],mul_res1[1167],mul_res1[1168],mul_res1[1169],mul_res1[1170],mul_res1[1171],mul_res1[1172],mul_res1[1173],mul_res1[1174],mul_res1[1175],mul_res1[1176],mul_res1[1177],mul_res1[1178],mul_res1[1179],mul_res1[1180],mul_res1[1181],mul_res1[1182],mul_res1[1183],mul_res1[1184],mul_res1[1185],mul_res1[1186],mul_res1[1187],mul_res1[1188],mul_res1[1189],mul_res1[1190],mul_res1[1191],mul_res1[1192],mul_res1[1193],mul_res1[1194],mul_res1[1195],mul_res1[1196],mul_res1[1197],mul_res1[1198],mul_res1[1199],result_fc1[5]);


adder_200in adder_200in_mod_6(clk,rst,mul_res1[1200],mul_res1[1201],mul_res1[1202],mul_res1[1203],mul_res1[1204],mul_res1[1205],mul_res1[1206],mul_res1[1207],mul_res1[1208],mul_res1[1209],mul_res1[1210],mul_res1[1211],mul_res1[1212],mul_res1[1213],mul_res1[1214],mul_res1[1215],mul_res1[1216],mul_res1[1217],mul_res1[1218],mul_res1[1219],mul_res1[1220],mul_res1[1221],mul_res1[1222],mul_res1[1223],mul_res1[1224],mul_res1[1225],mul_res1[1226],mul_res1[1227],mul_res1[1228],mul_res1[1229],mul_res1[1230],mul_res1[1231],mul_res1[1232],mul_res1[1233],mul_res1[1234],mul_res1[1235],mul_res1[1236],mul_res1[1237],mul_res1[1238],mul_res1[1239],mul_res1[1240],mul_res1[1241],mul_res1[1242],mul_res1[1243],mul_res1[1244],mul_res1[1245],mul_res1[1246],mul_res1[1247],mul_res1[1248],mul_res1[1249],mul_res1[1250],mul_res1[1251],mul_res1[1252],mul_res1[1253],mul_res1[1254],mul_res1[1255],mul_res1[1256],mul_res1[1257],mul_res1[1258],mul_res1[1259],mul_res1[1260],mul_res1[1261],mul_res1[1262],mul_res1[1263],mul_res1[1264],mul_res1[1265],mul_res1[1266],mul_res1[1267],mul_res1[1268],mul_res1[1269],mul_res1[1270],mul_res1[1271],mul_res1[1272],mul_res1[1273],mul_res1[1274],mul_res1[1275],mul_res1[1276],mul_res1[1277],mul_res1[1278],mul_res1[1279],mul_res1[1280],mul_res1[1281],mul_res1[1282],mul_res1[1283],mul_res1[1284],mul_res1[1285],mul_res1[1286],mul_res1[1287],mul_res1[1288],mul_res1[1289],mul_res1[1290],mul_res1[1291],mul_res1[1292],mul_res1[1293],mul_res1[1294],mul_res1[1295],mul_res1[1296],mul_res1[1297],mul_res1[1298],mul_res1[1299],mul_res1[1300],mul_res1[1301],mul_res1[1302],mul_res1[1303],mul_res1[1304],mul_res1[1305],mul_res1[1306],mul_res1[1307],mul_res1[1308],mul_res1[1309],mul_res1[1310],mul_res1[1311],mul_res1[1312],mul_res1[1313],mul_res1[1314],mul_res1[1315],mul_res1[1316],mul_res1[1317],mul_res1[1318],mul_res1[1319],mul_res1[1320],mul_res1[1321],mul_res1[1322],mul_res1[1323],mul_res1[1324],mul_res1[1325],mul_res1[1326],mul_res1[1327],mul_res1[1328],mul_res1[1329],mul_res1[1330],mul_res1[1331],mul_res1[1332],mul_res1[1333],mul_res1[1334],mul_res1[1335],mul_res1[1336],mul_res1[1337],mul_res1[1338],mul_res1[1339],mul_res1[1340],mul_res1[1341],mul_res1[1342],mul_res1[1343],mul_res1[1344],mul_res1[1345],mul_res1[1346],mul_res1[1347],mul_res1[1348],mul_res1[1349],mul_res1[1350],mul_res1[1351],mul_res1[1352],mul_res1[1353],mul_res1[1354],mul_res1[1355],mul_res1[1356],mul_res1[1357],mul_res1[1358],mul_res1[1359],mul_res1[1360],mul_res1[1361],mul_res1[1362],mul_res1[1363],mul_res1[1364],mul_res1[1365],mul_res1[1366],mul_res1[1367],mul_res1[1368],mul_res1[1369],mul_res1[1370],mul_res1[1371],mul_res1[1372],mul_res1[1373],mul_res1[1374],mul_res1[1375],mul_res1[1376],mul_res1[1377],mul_res1[1378],mul_res1[1379],mul_res1[1380],mul_res1[1381],mul_res1[1382],mul_res1[1383],mul_res1[1384],mul_res1[1385],mul_res1[1386],mul_res1[1387],mul_res1[1388],mul_res1[1389],mul_res1[1390],mul_res1[1391],mul_res1[1392],mul_res1[1393],mul_res1[1394],mul_res1[1395],mul_res1[1396],mul_res1[1397],mul_res1[1398],mul_res1[1399],result_fc1[6]);


adder_200in adder_200in_mod_7(clk,rst,mul_res1[1400],mul_res1[1401],mul_res1[1402],mul_res1[1403],mul_res1[1404],mul_res1[1405],mul_res1[1406],mul_res1[1407],mul_res1[1408],mul_res1[1409],mul_res1[1410],mul_res1[1411],mul_res1[1412],mul_res1[1413],mul_res1[1414],mul_res1[1415],mul_res1[1416],mul_res1[1417],mul_res1[1418],mul_res1[1419],mul_res1[1420],mul_res1[1421],mul_res1[1422],mul_res1[1423],mul_res1[1424],mul_res1[1425],mul_res1[1426],mul_res1[1427],mul_res1[1428],mul_res1[1429],mul_res1[1430],mul_res1[1431],mul_res1[1432],mul_res1[1433],mul_res1[1434],mul_res1[1435],mul_res1[1436],mul_res1[1437],mul_res1[1438],mul_res1[1439],mul_res1[1440],mul_res1[1441],mul_res1[1442],mul_res1[1443],mul_res1[1444],mul_res1[1445],mul_res1[1446],mul_res1[1447],mul_res1[1448],mul_res1[1449],mul_res1[1450],mul_res1[1451],mul_res1[1452],mul_res1[1453],mul_res1[1454],mul_res1[1455],mul_res1[1456],mul_res1[1457],mul_res1[1458],mul_res1[1459],mul_res1[1460],mul_res1[1461],mul_res1[1462],mul_res1[1463],mul_res1[1464],mul_res1[1465],mul_res1[1466],mul_res1[1467],mul_res1[1468],mul_res1[1469],mul_res1[1470],mul_res1[1471],mul_res1[1472],mul_res1[1473],mul_res1[1474],mul_res1[1475],mul_res1[1476],mul_res1[1477],mul_res1[1478],mul_res1[1479],mul_res1[1480],mul_res1[1481],mul_res1[1482],mul_res1[1483],mul_res1[1484],mul_res1[1485],mul_res1[1486],mul_res1[1487],mul_res1[1488],mul_res1[1489],mul_res1[1490],mul_res1[1491],mul_res1[1492],mul_res1[1493],mul_res1[1494],mul_res1[1495],mul_res1[1496],mul_res1[1497],mul_res1[1498],mul_res1[1499],mul_res1[1500],mul_res1[1501],mul_res1[1502],mul_res1[1503],mul_res1[1504],mul_res1[1505],mul_res1[1506],mul_res1[1507],mul_res1[1508],mul_res1[1509],mul_res1[1510],mul_res1[1511],mul_res1[1512],mul_res1[1513],mul_res1[1514],mul_res1[1515],mul_res1[1516],mul_res1[1517],mul_res1[1518],mul_res1[1519],mul_res1[1520],mul_res1[1521],mul_res1[1522],mul_res1[1523],mul_res1[1524],mul_res1[1525],mul_res1[1526],mul_res1[1527],mul_res1[1528],mul_res1[1529],mul_res1[1530],mul_res1[1531],mul_res1[1532],mul_res1[1533],mul_res1[1534],mul_res1[1535],mul_res1[1536],mul_res1[1537],mul_res1[1538],mul_res1[1539],mul_res1[1540],mul_res1[1541],mul_res1[1542],mul_res1[1543],mul_res1[1544],mul_res1[1545],mul_res1[1546],mul_res1[1547],mul_res1[1548],mul_res1[1549],mul_res1[1550],mul_res1[1551],mul_res1[1552],mul_res1[1553],mul_res1[1554],mul_res1[1555],mul_res1[1556],mul_res1[1557],mul_res1[1558],mul_res1[1559],mul_res1[1560],mul_res1[1561],mul_res1[1562],mul_res1[1563],mul_res1[1564],mul_res1[1565],mul_res1[1566],mul_res1[1567],mul_res1[1568],mul_res1[1569],mul_res1[1570],mul_res1[1571],mul_res1[1572],mul_res1[1573],mul_res1[1574],mul_res1[1575],mul_res1[1576],mul_res1[1577],mul_res1[1578],mul_res1[1579],mul_res1[1580],mul_res1[1581],mul_res1[1582],mul_res1[1583],mul_res1[1584],mul_res1[1585],mul_res1[1586],mul_res1[1587],mul_res1[1588],mul_res1[1589],mul_res1[1590],mul_res1[1591],mul_res1[1592],mul_res1[1593],mul_res1[1594],mul_res1[1595],mul_res1[1596],mul_res1[1597],mul_res1[1598],mul_res1[1599],result_fc1[7]);


adder_200in adder_200in_mod_8(clk,rst,mul_res1[1600],mul_res1[1601],mul_res1[1602],mul_res1[1603],mul_res1[1604],mul_res1[1605],mul_res1[1606],mul_res1[1607],mul_res1[1608],mul_res1[1609],mul_res1[1610],mul_res1[1611],mul_res1[1612],mul_res1[1613],mul_res1[1614],mul_res1[1615],mul_res1[1616],mul_res1[1617],mul_res1[1618],mul_res1[1619],mul_res1[1620],mul_res1[1621],mul_res1[1622],mul_res1[1623],mul_res1[1624],mul_res1[1625],mul_res1[1626],mul_res1[1627],mul_res1[1628],mul_res1[1629],mul_res1[1630],mul_res1[1631],mul_res1[1632],mul_res1[1633],mul_res1[1634],mul_res1[1635],mul_res1[1636],mul_res1[1637],mul_res1[1638],mul_res1[1639],mul_res1[1640],mul_res1[1641],mul_res1[1642],mul_res1[1643],mul_res1[1644],mul_res1[1645],mul_res1[1646],mul_res1[1647],mul_res1[1648],mul_res1[1649],mul_res1[1650],mul_res1[1651],mul_res1[1652],mul_res1[1653],mul_res1[1654],mul_res1[1655],mul_res1[1656],mul_res1[1657],mul_res1[1658],mul_res1[1659],mul_res1[1660],mul_res1[1661],mul_res1[1662],mul_res1[1663],mul_res1[1664],mul_res1[1665],mul_res1[1666],mul_res1[1667],mul_res1[1668],mul_res1[1669],mul_res1[1670],mul_res1[1671],mul_res1[1672],mul_res1[1673],mul_res1[1674],mul_res1[1675],mul_res1[1676],mul_res1[1677],mul_res1[1678],mul_res1[1679],mul_res1[1680],mul_res1[1681],mul_res1[1682],mul_res1[1683],mul_res1[1684],mul_res1[1685],mul_res1[1686],mul_res1[1687],mul_res1[1688],mul_res1[1689],mul_res1[1690],mul_res1[1691],mul_res1[1692],mul_res1[1693],mul_res1[1694],mul_res1[1695],mul_res1[1696],mul_res1[1697],mul_res1[1698],mul_res1[1699],mul_res1[1700],mul_res1[1701],mul_res1[1702],mul_res1[1703],mul_res1[1704],mul_res1[1705],mul_res1[1706],mul_res1[1707],mul_res1[1708],mul_res1[1709],mul_res1[1710],mul_res1[1711],mul_res1[1712],mul_res1[1713],mul_res1[1714],mul_res1[1715],mul_res1[1716],mul_res1[1717],mul_res1[1718],mul_res1[1719],mul_res1[1720],mul_res1[1721],mul_res1[1722],mul_res1[1723],mul_res1[1724],mul_res1[1725],mul_res1[1726],mul_res1[1727],mul_res1[1728],mul_res1[1729],mul_res1[1730],mul_res1[1731],mul_res1[1732],mul_res1[1733],mul_res1[1734],mul_res1[1735],mul_res1[1736],mul_res1[1737],mul_res1[1738],mul_res1[1739],mul_res1[1740],mul_res1[1741],mul_res1[1742],mul_res1[1743],mul_res1[1744],mul_res1[1745],mul_res1[1746],mul_res1[1747],mul_res1[1748],mul_res1[1749],mul_res1[1750],mul_res1[1751],mul_res1[1752],mul_res1[1753],mul_res1[1754],mul_res1[1755],mul_res1[1756],mul_res1[1757],mul_res1[1758],mul_res1[1759],mul_res1[1760],mul_res1[1761],mul_res1[1762],mul_res1[1763],mul_res1[1764],mul_res1[1765],mul_res1[1766],mul_res1[1767],mul_res1[1768],mul_res1[1769],mul_res1[1770],mul_res1[1771],mul_res1[1772],mul_res1[1773],mul_res1[1774],mul_res1[1775],mul_res1[1776],mul_res1[1777],mul_res1[1778],mul_res1[1779],mul_res1[1780],mul_res1[1781],mul_res1[1782],mul_res1[1783],mul_res1[1784],mul_res1[1785],mul_res1[1786],mul_res1[1787],mul_res1[1788],mul_res1[1789],mul_res1[1790],mul_res1[1791],mul_res1[1792],mul_res1[1793],mul_res1[1794],mul_res1[1795],mul_res1[1796],mul_res1[1797],mul_res1[1798],mul_res1[1799],result_fc1[8]);


adder_200in adder_200in_mod_9(clk,rst,mul_res1[1800],mul_res1[1801],mul_res1[1802],mul_res1[1803],mul_res1[1804],mul_res1[1805],mul_res1[1806],mul_res1[1807],mul_res1[1808],mul_res1[1809],mul_res1[1810],mul_res1[1811],mul_res1[1812],mul_res1[1813],mul_res1[1814],mul_res1[1815],mul_res1[1816],mul_res1[1817],mul_res1[1818],mul_res1[1819],mul_res1[1820],mul_res1[1821],mul_res1[1822],mul_res1[1823],mul_res1[1824],mul_res1[1825],mul_res1[1826],mul_res1[1827],mul_res1[1828],mul_res1[1829],mul_res1[1830],mul_res1[1831],mul_res1[1832],mul_res1[1833],mul_res1[1834],mul_res1[1835],mul_res1[1836],mul_res1[1837],mul_res1[1838],mul_res1[1839],mul_res1[1840],mul_res1[1841],mul_res1[1842],mul_res1[1843],mul_res1[1844],mul_res1[1845],mul_res1[1846],mul_res1[1847],mul_res1[1848],mul_res1[1849],mul_res1[1850],mul_res1[1851],mul_res1[1852],mul_res1[1853],mul_res1[1854],mul_res1[1855],mul_res1[1856],mul_res1[1857],mul_res1[1858],mul_res1[1859],mul_res1[1860],mul_res1[1861],mul_res1[1862],mul_res1[1863],mul_res1[1864],mul_res1[1865],mul_res1[1866],mul_res1[1867],mul_res1[1868],mul_res1[1869],mul_res1[1870],mul_res1[1871],mul_res1[1872],mul_res1[1873],mul_res1[1874],mul_res1[1875],mul_res1[1876],mul_res1[1877],mul_res1[1878],mul_res1[1879],mul_res1[1880],mul_res1[1881],mul_res1[1882],mul_res1[1883],mul_res1[1884],mul_res1[1885],mul_res1[1886],mul_res1[1887],mul_res1[1888],mul_res1[1889],mul_res1[1890],mul_res1[1891],mul_res1[1892],mul_res1[1893],mul_res1[1894],mul_res1[1895],mul_res1[1896],mul_res1[1897],mul_res1[1898],mul_res1[1899],mul_res1[1900],mul_res1[1901],mul_res1[1902],mul_res1[1903],mul_res1[1904],mul_res1[1905],mul_res1[1906],mul_res1[1907],mul_res1[1908],mul_res1[1909],mul_res1[1910],mul_res1[1911],mul_res1[1912],mul_res1[1913],mul_res1[1914],mul_res1[1915],mul_res1[1916],mul_res1[1917],mul_res1[1918],mul_res1[1919],mul_res1[1920],mul_res1[1921],mul_res1[1922],mul_res1[1923],mul_res1[1924],mul_res1[1925],mul_res1[1926],mul_res1[1927],mul_res1[1928],mul_res1[1929],mul_res1[1930],mul_res1[1931],mul_res1[1932],mul_res1[1933],mul_res1[1934],mul_res1[1935],mul_res1[1936],mul_res1[1937],mul_res1[1938],mul_res1[1939],mul_res1[1940],mul_res1[1941],mul_res1[1942],mul_res1[1943],mul_res1[1944],mul_res1[1945],mul_res1[1946],mul_res1[1947],mul_res1[1948],mul_res1[1949],mul_res1[1950],mul_res1[1951],mul_res1[1952],mul_res1[1953],mul_res1[1954],mul_res1[1955],mul_res1[1956],mul_res1[1957],mul_res1[1958],mul_res1[1959],mul_res1[1960],mul_res1[1961],mul_res1[1962],mul_res1[1963],mul_res1[1964],mul_res1[1965],mul_res1[1966],mul_res1[1967],mul_res1[1968],mul_res1[1969],mul_res1[1970],mul_res1[1971],mul_res1[1972],mul_res1[1973],mul_res1[1974],mul_res1[1975],mul_res1[1976],mul_res1[1977],mul_res1[1978],mul_res1[1979],mul_res1[1980],mul_res1[1981],mul_res1[1982],mul_res1[1983],mul_res1[1984],mul_res1[1985],mul_res1[1986],mul_res1[1987],mul_res1[1988],mul_res1[1989],mul_res1[1990],mul_res1[1991],mul_res1[1992],mul_res1[1993],mul_res1[1994],mul_res1[1995],mul_res1[1996],mul_res1[1997],mul_res1[1998],mul_res1[1999],result_fc1[9]);


adder_200in adder_200in_mod_10(clk,rst,mul_res1[2000],mul_res1[2001],mul_res1[2002],mul_res1[2003],mul_res1[2004],mul_res1[2005],mul_res1[2006],mul_res1[2007],mul_res1[2008],mul_res1[2009],mul_res1[2010],mul_res1[2011],mul_res1[2012],mul_res1[2013],mul_res1[2014],mul_res1[2015],mul_res1[2016],mul_res1[2017],mul_res1[2018],mul_res1[2019],mul_res1[2020],mul_res1[2021],mul_res1[2022],mul_res1[2023],mul_res1[2024],mul_res1[2025],mul_res1[2026],mul_res1[2027],mul_res1[2028],mul_res1[2029],mul_res1[2030],mul_res1[2031],mul_res1[2032],mul_res1[2033],mul_res1[2034],mul_res1[2035],mul_res1[2036],mul_res1[2037],mul_res1[2038],mul_res1[2039],mul_res1[2040],mul_res1[2041],mul_res1[2042],mul_res1[2043],mul_res1[2044],mul_res1[2045],mul_res1[2046],mul_res1[2047],mul_res1[2048],mul_res1[2049],mul_res1[2050],mul_res1[2051],mul_res1[2052],mul_res1[2053],mul_res1[2054],mul_res1[2055],mul_res1[2056],mul_res1[2057],mul_res1[2058],mul_res1[2059],mul_res1[2060],mul_res1[2061],mul_res1[2062],mul_res1[2063],mul_res1[2064],mul_res1[2065],mul_res1[2066],mul_res1[2067],mul_res1[2068],mul_res1[2069],mul_res1[2070],mul_res1[2071],mul_res1[2072],mul_res1[2073],mul_res1[2074],mul_res1[2075],mul_res1[2076],mul_res1[2077],mul_res1[2078],mul_res1[2079],mul_res1[2080],mul_res1[2081],mul_res1[2082],mul_res1[2083],mul_res1[2084],mul_res1[2085],mul_res1[2086],mul_res1[2087],mul_res1[2088],mul_res1[2089],mul_res1[2090],mul_res1[2091],mul_res1[2092],mul_res1[2093],mul_res1[2094],mul_res1[2095],mul_res1[2096],mul_res1[2097],mul_res1[2098],mul_res1[2099],mul_res1[2100],mul_res1[2101],mul_res1[2102],mul_res1[2103],mul_res1[2104],mul_res1[2105],mul_res1[2106],mul_res1[2107],mul_res1[2108],mul_res1[2109],mul_res1[2110],mul_res1[2111],mul_res1[2112],mul_res1[2113],mul_res1[2114],mul_res1[2115],mul_res1[2116],mul_res1[2117],mul_res1[2118],mul_res1[2119],mul_res1[2120],mul_res1[2121],mul_res1[2122],mul_res1[2123],mul_res1[2124],mul_res1[2125],mul_res1[2126],mul_res1[2127],mul_res1[2128],mul_res1[2129],mul_res1[2130],mul_res1[2131],mul_res1[2132],mul_res1[2133],mul_res1[2134],mul_res1[2135],mul_res1[2136],mul_res1[2137],mul_res1[2138],mul_res1[2139],mul_res1[2140],mul_res1[2141],mul_res1[2142],mul_res1[2143],mul_res1[2144],mul_res1[2145],mul_res1[2146],mul_res1[2147],mul_res1[2148],mul_res1[2149],mul_res1[2150],mul_res1[2151],mul_res1[2152],mul_res1[2153],mul_res1[2154],mul_res1[2155],mul_res1[2156],mul_res1[2157],mul_res1[2158],mul_res1[2159],mul_res1[2160],mul_res1[2161],mul_res1[2162],mul_res1[2163],mul_res1[2164],mul_res1[2165],mul_res1[2166],mul_res1[2167],mul_res1[2168],mul_res1[2169],mul_res1[2170],mul_res1[2171],mul_res1[2172],mul_res1[2173],mul_res1[2174],mul_res1[2175],mul_res1[2176],mul_res1[2177],mul_res1[2178],mul_res1[2179],mul_res1[2180],mul_res1[2181],mul_res1[2182],mul_res1[2183],mul_res1[2184],mul_res1[2185],mul_res1[2186],mul_res1[2187],mul_res1[2188],mul_res1[2189],mul_res1[2190],mul_res1[2191],mul_res1[2192],mul_res1[2193],mul_res1[2194],mul_res1[2195],mul_res1[2196],mul_res1[2197],mul_res1[2198],mul_res1[2199],result_fc1[10]);


adder_200in adder_200in_mod_11(clk,rst,mul_res1[2200],mul_res1[2201],mul_res1[2202],mul_res1[2203],mul_res1[2204],mul_res1[2205],mul_res1[2206],mul_res1[2207],mul_res1[2208],mul_res1[2209],mul_res1[2210],mul_res1[2211],mul_res1[2212],mul_res1[2213],mul_res1[2214],mul_res1[2215],mul_res1[2216],mul_res1[2217],mul_res1[2218],mul_res1[2219],mul_res1[2220],mul_res1[2221],mul_res1[2222],mul_res1[2223],mul_res1[2224],mul_res1[2225],mul_res1[2226],mul_res1[2227],mul_res1[2228],mul_res1[2229],mul_res1[2230],mul_res1[2231],mul_res1[2232],mul_res1[2233],mul_res1[2234],mul_res1[2235],mul_res1[2236],mul_res1[2237],mul_res1[2238],mul_res1[2239],mul_res1[2240],mul_res1[2241],mul_res1[2242],mul_res1[2243],mul_res1[2244],mul_res1[2245],mul_res1[2246],mul_res1[2247],mul_res1[2248],mul_res1[2249],mul_res1[2250],mul_res1[2251],mul_res1[2252],mul_res1[2253],mul_res1[2254],mul_res1[2255],mul_res1[2256],mul_res1[2257],mul_res1[2258],mul_res1[2259],mul_res1[2260],mul_res1[2261],mul_res1[2262],mul_res1[2263],mul_res1[2264],mul_res1[2265],mul_res1[2266],mul_res1[2267],mul_res1[2268],mul_res1[2269],mul_res1[2270],mul_res1[2271],mul_res1[2272],mul_res1[2273],mul_res1[2274],mul_res1[2275],mul_res1[2276],mul_res1[2277],mul_res1[2278],mul_res1[2279],mul_res1[2280],mul_res1[2281],mul_res1[2282],mul_res1[2283],mul_res1[2284],mul_res1[2285],mul_res1[2286],mul_res1[2287],mul_res1[2288],mul_res1[2289],mul_res1[2290],mul_res1[2291],mul_res1[2292],mul_res1[2293],mul_res1[2294],mul_res1[2295],mul_res1[2296],mul_res1[2297],mul_res1[2298],mul_res1[2299],mul_res1[2300],mul_res1[2301],mul_res1[2302],mul_res1[2303],mul_res1[2304],mul_res1[2305],mul_res1[2306],mul_res1[2307],mul_res1[2308],mul_res1[2309],mul_res1[2310],mul_res1[2311],mul_res1[2312],mul_res1[2313],mul_res1[2314],mul_res1[2315],mul_res1[2316],mul_res1[2317],mul_res1[2318],mul_res1[2319],mul_res1[2320],mul_res1[2321],mul_res1[2322],mul_res1[2323],mul_res1[2324],mul_res1[2325],mul_res1[2326],mul_res1[2327],mul_res1[2328],mul_res1[2329],mul_res1[2330],mul_res1[2331],mul_res1[2332],mul_res1[2333],mul_res1[2334],mul_res1[2335],mul_res1[2336],mul_res1[2337],mul_res1[2338],mul_res1[2339],mul_res1[2340],mul_res1[2341],mul_res1[2342],mul_res1[2343],mul_res1[2344],mul_res1[2345],mul_res1[2346],mul_res1[2347],mul_res1[2348],mul_res1[2349],mul_res1[2350],mul_res1[2351],mul_res1[2352],mul_res1[2353],mul_res1[2354],mul_res1[2355],mul_res1[2356],mul_res1[2357],mul_res1[2358],mul_res1[2359],mul_res1[2360],mul_res1[2361],mul_res1[2362],mul_res1[2363],mul_res1[2364],mul_res1[2365],mul_res1[2366],mul_res1[2367],mul_res1[2368],mul_res1[2369],mul_res1[2370],mul_res1[2371],mul_res1[2372],mul_res1[2373],mul_res1[2374],mul_res1[2375],mul_res1[2376],mul_res1[2377],mul_res1[2378],mul_res1[2379],mul_res1[2380],mul_res1[2381],mul_res1[2382],mul_res1[2383],mul_res1[2384],mul_res1[2385],mul_res1[2386],mul_res1[2387],mul_res1[2388],mul_res1[2389],mul_res1[2390],mul_res1[2391],mul_res1[2392],mul_res1[2393],mul_res1[2394],mul_res1[2395],mul_res1[2396],mul_res1[2397],mul_res1[2398],mul_res1[2399],result_fc1[11]);


adder_200in adder_200in_mod_12(clk,rst,mul_res1[2400],mul_res1[2401],mul_res1[2402],mul_res1[2403],mul_res1[2404],mul_res1[2405],mul_res1[2406],mul_res1[2407],mul_res1[2408],mul_res1[2409],mul_res1[2410],mul_res1[2411],mul_res1[2412],mul_res1[2413],mul_res1[2414],mul_res1[2415],mul_res1[2416],mul_res1[2417],mul_res1[2418],mul_res1[2419],mul_res1[2420],mul_res1[2421],mul_res1[2422],mul_res1[2423],mul_res1[2424],mul_res1[2425],mul_res1[2426],mul_res1[2427],mul_res1[2428],mul_res1[2429],mul_res1[2430],mul_res1[2431],mul_res1[2432],mul_res1[2433],mul_res1[2434],mul_res1[2435],mul_res1[2436],mul_res1[2437],mul_res1[2438],mul_res1[2439],mul_res1[2440],mul_res1[2441],mul_res1[2442],mul_res1[2443],mul_res1[2444],mul_res1[2445],mul_res1[2446],mul_res1[2447],mul_res1[2448],mul_res1[2449],mul_res1[2450],mul_res1[2451],mul_res1[2452],mul_res1[2453],mul_res1[2454],mul_res1[2455],mul_res1[2456],mul_res1[2457],mul_res1[2458],mul_res1[2459],mul_res1[2460],mul_res1[2461],mul_res1[2462],mul_res1[2463],mul_res1[2464],mul_res1[2465],mul_res1[2466],mul_res1[2467],mul_res1[2468],mul_res1[2469],mul_res1[2470],mul_res1[2471],mul_res1[2472],mul_res1[2473],mul_res1[2474],mul_res1[2475],mul_res1[2476],mul_res1[2477],mul_res1[2478],mul_res1[2479],mul_res1[2480],mul_res1[2481],mul_res1[2482],mul_res1[2483],mul_res1[2484],mul_res1[2485],mul_res1[2486],mul_res1[2487],mul_res1[2488],mul_res1[2489],mul_res1[2490],mul_res1[2491],mul_res1[2492],mul_res1[2493],mul_res1[2494],mul_res1[2495],mul_res1[2496],mul_res1[2497],mul_res1[2498],mul_res1[2499],mul_res1[2500],mul_res1[2501],mul_res1[2502],mul_res1[2503],mul_res1[2504],mul_res1[2505],mul_res1[2506],mul_res1[2507],mul_res1[2508],mul_res1[2509],mul_res1[2510],mul_res1[2511],mul_res1[2512],mul_res1[2513],mul_res1[2514],mul_res1[2515],mul_res1[2516],mul_res1[2517],mul_res1[2518],mul_res1[2519],mul_res1[2520],mul_res1[2521],mul_res1[2522],mul_res1[2523],mul_res1[2524],mul_res1[2525],mul_res1[2526],mul_res1[2527],mul_res1[2528],mul_res1[2529],mul_res1[2530],mul_res1[2531],mul_res1[2532],mul_res1[2533],mul_res1[2534],mul_res1[2535],mul_res1[2536],mul_res1[2537],mul_res1[2538],mul_res1[2539],mul_res1[2540],mul_res1[2541],mul_res1[2542],mul_res1[2543],mul_res1[2544],mul_res1[2545],mul_res1[2546],mul_res1[2547],mul_res1[2548],mul_res1[2549],mul_res1[2550],mul_res1[2551],mul_res1[2552],mul_res1[2553],mul_res1[2554],mul_res1[2555],mul_res1[2556],mul_res1[2557],mul_res1[2558],mul_res1[2559],mul_res1[2560],mul_res1[2561],mul_res1[2562],mul_res1[2563],mul_res1[2564],mul_res1[2565],mul_res1[2566],mul_res1[2567],mul_res1[2568],mul_res1[2569],mul_res1[2570],mul_res1[2571],mul_res1[2572],mul_res1[2573],mul_res1[2574],mul_res1[2575],mul_res1[2576],mul_res1[2577],mul_res1[2578],mul_res1[2579],mul_res1[2580],mul_res1[2581],mul_res1[2582],mul_res1[2583],mul_res1[2584],mul_res1[2585],mul_res1[2586],mul_res1[2587],mul_res1[2588],mul_res1[2589],mul_res1[2590],mul_res1[2591],mul_res1[2592],mul_res1[2593],mul_res1[2594],mul_res1[2595],mul_res1[2596],mul_res1[2597],mul_res1[2598],mul_res1[2599],result_fc1[12]);


adder_200in adder_200in_mod_13(clk,rst,mul_res1[2600],mul_res1[2601],mul_res1[2602],mul_res1[2603],mul_res1[2604],mul_res1[2605],mul_res1[2606],mul_res1[2607],mul_res1[2608],mul_res1[2609],mul_res1[2610],mul_res1[2611],mul_res1[2612],mul_res1[2613],mul_res1[2614],mul_res1[2615],mul_res1[2616],mul_res1[2617],mul_res1[2618],mul_res1[2619],mul_res1[2620],mul_res1[2621],mul_res1[2622],mul_res1[2623],mul_res1[2624],mul_res1[2625],mul_res1[2626],mul_res1[2627],mul_res1[2628],mul_res1[2629],mul_res1[2630],mul_res1[2631],mul_res1[2632],mul_res1[2633],mul_res1[2634],mul_res1[2635],mul_res1[2636],mul_res1[2637],mul_res1[2638],mul_res1[2639],mul_res1[2640],mul_res1[2641],mul_res1[2642],mul_res1[2643],mul_res1[2644],mul_res1[2645],mul_res1[2646],mul_res1[2647],mul_res1[2648],mul_res1[2649],mul_res1[2650],mul_res1[2651],mul_res1[2652],mul_res1[2653],mul_res1[2654],mul_res1[2655],mul_res1[2656],mul_res1[2657],mul_res1[2658],mul_res1[2659],mul_res1[2660],mul_res1[2661],mul_res1[2662],mul_res1[2663],mul_res1[2664],mul_res1[2665],mul_res1[2666],mul_res1[2667],mul_res1[2668],mul_res1[2669],mul_res1[2670],mul_res1[2671],mul_res1[2672],mul_res1[2673],mul_res1[2674],mul_res1[2675],mul_res1[2676],mul_res1[2677],mul_res1[2678],mul_res1[2679],mul_res1[2680],mul_res1[2681],mul_res1[2682],mul_res1[2683],mul_res1[2684],mul_res1[2685],mul_res1[2686],mul_res1[2687],mul_res1[2688],mul_res1[2689],mul_res1[2690],mul_res1[2691],mul_res1[2692],mul_res1[2693],mul_res1[2694],mul_res1[2695],mul_res1[2696],mul_res1[2697],mul_res1[2698],mul_res1[2699],mul_res1[2700],mul_res1[2701],mul_res1[2702],mul_res1[2703],mul_res1[2704],mul_res1[2705],mul_res1[2706],mul_res1[2707],mul_res1[2708],mul_res1[2709],mul_res1[2710],mul_res1[2711],mul_res1[2712],mul_res1[2713],mul_res1[2714],mul_res1[2715],mul_res1[2716],mul_res1[2717],mul_res1[2718],mul_res1[2719],mul_res1[2720],mul_res1[2721],mul_res1[2722],mul_res1[2723],mul_res1[2724],mul_res1[2725],mul_res1[2726],mul_res1[2727],mul_res1[2728],mul_res1[2729],mul_res1[2730],mul_res1[2731],mul_res1[2732],mul_res1[2733],mul_res1[2734],mul_res1[2735],mul_res1[2736],mul_res1[2737],mul_res1[2738],mul_res1[2739],mul_res1[2740],mul_res1[2741],mul_res1[2742],mul_res1[2743],mul_res1[2744],mul_res1[2745],mul_res1[2746],mul_res1[2747],mul_res1[2748],mul_res1[2749],mul_res1[2750],mul_res1[2751],mul_res1[2752],mul_res1[2753],mul_res1[2754],mul_res1[2755],mul_res1[2756],mul_res1[2757],mul_res1[2758],mul_res1[2759],mul_res1[2760],mul_res1[2761],mul_res1[2762],mul_res1[2763],mul_res1[2764],mul_res1[2765],mul_res1[2766],mul_res1[2767],mul_res1[2768],mul_res1[2769],mul_res1[2770],mul_res1[2771],mul_res1[2772],mul_res1[2773],mul_res1[2774],mul_res1[2775],mul_res1[2776],mul_res1[2777],mul_res1[2778],mul_res1[2779],mul_res1[2780],mul_res1[2781],mul_res1[2782],mul_res1[2783],mul_res1[2784],mul_res1[2785],mul_res1[2786],mul_res1[2787],mul_res1[2788],mul_res1[2789],mul_res1[2790],mul_res1[2791],mul_res1[2792],mul_res1[2793],mul_res1[2794],mul_res1[2795],mul_res1[2796],mul_res1[2797],mul_res1[2798],mul_res1[2799],result_fc1[13]);


adder_200in adder_200in_mod_14(clk,rst,mul_res1[2800],mul_res1[2801],mul_res1[2802],mul_res1[2803],mul_res1[2804],mul_res1[2805],mul_res1[2806],mul_res1[2807],mul_res1[2808],mul_res1[2809],mul_res1[2810],mul_res1[2811],mul_res1[2812],mul_res1[2813],mul_res1[2814],mul_res1[2815],mul_res1[2816],mul_res1[2817],mul_res1[2818],mul_res1[2819],mul_res1[2820],mul_res1[2821],mul_res1[2822],mul_res1[2823],mul_res1[2824],mul_res1[2825],mul_res1[2826],mul_res1[2827],mul_res1[2828],mul_res1[2829],mul_res1[2830],mul_res1[2831],mul_res1[2832],mul_res1[2833],mul_res1[2834],mul_res1[2835],mul_res1[2836],mul_res1[2837],mul_res1[2838],mul_res1[2839],mul_res1[2840],mul_res1[2841],mul_res1[2842],mul_res1[2843],mul_res1[2844],mul_res1[2845],mul_res1[2846],mul_res1[2847],mul_res1[2848],mul_res1[2849],mul_res1[2850],mul_res1[2851],mul_res1[2852],mul_res1[2853],mul_res1[2854],mul_res1[2855],mul_res1[2856],mul_res1[2857],mul_res1[2858],mul_res1[2859],mul_res1[2860],mul_res1[2861],mul_res1[2862],mul_res1[2863],mul_res1[2864],mul_res1[2865],mul_res1[2866],mul_res1[2867],mul_res1[2868],mul_res1[2869],mul_res1[2870],mul_res1[2871],mul_res1[2872],mul_res1[2873],mul_res1[2874],mul_res1[2875],mul_res1[2876],mul_res1[2877],mul_res1[2878],mul_res1[2879],mul_res1[2880],mul_res1[2881],mul_res1[2882],mul_res1[2883],mul_res1[2884],mul_res1[2885],mul_res1[2886],mul_res1[2887],mul_res1[2888],mul_res1[2889],mul_res1[2890],mul_res1[2891],mul_res1[2892],mul_res1[2893],mul_res1[2894],mul_res1[2895],mul_res1[2896],mul_res1[2897],mul_res1[2898],mul_res1[2899],mul_res1[2900],mul_res1[2901],mul_res1[2902],mul_res1[2903],mul_res1[2904],mul_res1[2905],mul_res1[2906],mul_res1[2907],mul_res1[2908],mul_res1[2909],mul_res1[2910],mul_res1[2911],mul_res1[2912],mul_res1[2913],mul_res1[2914],mul_res1[2915],mul_res1[2916],mul_res1[2917],mul_res1[2918],mul_res1[2919],mul_res1[2920],mul_res1[2921],mul_res1[2922],mul_res1[2923],mul_res1[2924],mul_res1[2925],mul_res1[2926],mul_res1[2927],mul_res1[2928],mul_res1[2929],mul_res1[2930],mul_res1[2931],mul_res1[2932],mul_res1[2933],mul_res1[2934],mul_res1[2935],mul_res1[2936],mul_res1[2937],mul_res1[2938],mul_res1[2939],mul_res1[2940],mul_res1[2941],mul_res1[2942],mul_res1[2943],mul_res1[2944],mul_res1[2945],mul_res1[2946],mul_res1[2947],mul_res1[2948],mul_res1[2949],mul_res1[2950],mul_res1[2951],mul_res1[2952],mul_res1[2953],mul_res1[2954],mul_res1[2955],mul_res1[2956],mul_res1[2957],mul_res1[2958],mul_res1[2959],mul_res1[2960],mul_res1[2961],mul_res1[2962],mul_res1[2963],mul_res1[2964],mul_res1[2965],mul_res1[2966],mul_res1[2967],mul_res1[2968],mul_res1[2969],mul_res1[2970],mul_res1[2971],mul_res1[2972],mul_res1[2973],mul_res1[2974],mul_res1[2975],mul_res1[2976],mul_res1[2977],mul_res1[2978],mul_res1[2979],mul_res1[2980],mul_res1[2981],mul_res1[2982],mul_res1[2983],mul_res1[2984],mul_res1[2985],mul_res1[2986],mul_res1[2987],mul_res1[2988],mul_res1[2989],mul_res1[2990],mul_res1[2991],mul_res1[2992],mul_res1[2993],mul_res1[2994],mul_res1[2995],mul_res1[2996],mul_res1[2997],mul_res1[2998],mul_res1[2999],result_fc1[14]);


adder_200in adder_200in_mod_15(clk,rst,mul_res1[3000],mul_res1[3001],mul_res1[3002],mul_res1[3003],mul_res1[3004],mul_res1[3005],mul_res1[3006],mul_res1[3007],mul_res1[3008],mul_res1[3009],mul_res1[3010],mul_res1[3011],mul_res1[3012],mul_res1[3013],mul_res1[3014],mul_res1[3015],mul_res1[3016],mul_res1[3017],mul_res1[3018],mul_res1[3019],mul_res1[3020],mul_res1[3021],mul_res1[3022],mul_res1[3023],mul_res1[3024],mul_res1[3025],mul_res1[3026],mul_res1[3027],mul_res1[3028],mul_res1[3029],mul_res1[3030],mul_res1[3031],mul_res1[3032],mul_res1[3033],mul_res1[3034],mul_res1[3035],mul_res1[3036],mul_res1[3037],mul_res1[3038],mul_res1[3039],mul_res1[3040],mul_res1[3041],mul_res1[3042],mul_res1[3043],mul_res1[3044],mul_res1[3045],mul_res1[3046],mul_res1[3047],mul_res1[3048],mul_res1[3049],mul_res1[3050],mul_res1[3051],mul_res1[3052],mul_res1[3053],mul_res1[3054],mul_res1[3055],mul_res1[3056],mul_res1[3057],mul_res1[3058],mul_res1[3059],mul_res1[3060],mul_res1[3061],mul_res1[3062],mul_res1[3063],mul_res1[3064],mul_res1[3065],mul_res1[3066],mul_res1[3067],mul_res1[3068],mul_res1[3069],mul_res1[3070],mul_res1[3071],mul_res1[3072],mul_res1[3073],mul_res1[3074],mul_res1[3075],mul_res1[3076],mul_res1[3077],mul_res1[3078],mul_res1[3079],mul_res1[3080],mul_res1[3081],mul_res1[3082],mul_res1[3083],mul_res1[3084],mul_res1[3085],mul_res1[3086],mul_res1[3087],mul_res1[3088],mul_res1[3089],mul_res1[3090],mul_res1[3091],mul_res1[3092],mul_res1[3093],mul_res1[3094],mul_res1[3095],mul_res1[3096],mul_res1[3097],mul_res1[3098],mul_res1[3099],mul_res1[3100],mul_res1[3101],mul_res1[3102],mul_res1[3103],mul_res1[3104],mul_res1[3105],mul_res1[3106],mul_res1[3107],mul_res1[3108],mul_res1[3109],mul_res1[3110],mul_res1[3111],mul_res1[3112],mul_res1[3113],mul_res1[3114],mul_res1[3115],mul_res1[3116],mul_res1[3117],mul_res1[3118],mul_res1[3119],mul_res1[3120],mul_res1[3121],mul_res1[3122],mul_res1[3123],mul_res1[3124],mul_res1[3125],mul_res1[3126],mul_res1[3127],mul_res1[3128],mul_res1[3129],mul_res1[3130],mul_res1[3131],mul_res1[3132],mul_res1[3133],mul_res1[3134],mul_res1[3135],mul_res1[3136],mul_res1[3137],mul_res1[3138],mul_res1[3139],mul_res1[3140],mul_res1[3141],mul_res1[3142],mul_res1[3143],mul_res1[3144],mul_res1[3145],mul_res1[3146],mul_res1[3147],mul_res1[3148],mul_res1[3149],mul_res1[3150],mul_res1[3151],mul_res1[3152],mul_res1[3153],mul_res1[3154],mul_res1[3155],mul_res1[3156],mul_res1[3157],mul_res1[3158],mul_res1[3159],mul_res1[3160],mul_res1[3161],mul_res1[3162],mul_res1[3163],mul_res1[3164],mul_res1[3165],mul_res1[3166],mul_res1[3167],mul_res1[3168],mul_res1[3169],mul_res1[3170],mul_res1[3171],mul_res1[3172],mul_res1[3173],mul_res1[3174],mul_res1[3175],mul_res1[3176],mul_res1[3177],mul_res1[3178],mul_res1[3179],mul_res1[3180],mul_res1[3181],mul_res1[3182],mul_res1[3183],mul_res1[3184],mul_res1[3185],mul_res1[3186],mul_res1[3187],mul_res1[3188],mul_res1[3189],mul_res1[3190],mul_res1[3191],mul_res1[3192],mul_res1[3193],mul_res1[3194],mul_res1[3195],mul_res1[3196],mul_res1[3197],mul_res1[3198],mul_res1[3199],result_fc1[15]);


adder_200in adder_200in_mod_16(clk,rst,mul_res1[3200],mul_res1[3201],mul_res1[3202],mul_res1[3203],mul_res1[3204],mul_res1[3205],mul_res1[3206],mul_res1[3207],mul_res1[3208],mul_res1[3209],mul_res1[3210],mul_res1[3211],mul_res1[3212],mul_res1[3213],mul_res1[3214],mul_res1[3215],mul_res1[3216],mul_res1[3217],mul_res1[3218],mul_res1[3219],mul_res1[3220],mul_res1[3221],mul_res1[3222],mul_res1[3223],mul_res1[3224],mul_res1[3225],mul_res1[3226],mul_res1[3227],mul_res1[3228],mul_res1[3229],mul_res1[3230],mul_res1[3231],mul_res1[3232],mul_res1[3233],mul_res1[3234],mul_res1[3235],mul_res1[3236],mul_res1[3237],mul_res1[3238],mul_res1[3239],mul_res1[3240],mul_res1[3241],mul_res1[3242],mul_res1[3243],mul_res1[3244],mul_res1[3245],mul_res1[3246],mul_res1[3247],mul_res1[3248],mul_res1[3249],mul_res1[3250],mul_res1[3251],mul_res1[3252],mul_res1[3253],mul_res1[3254],mul_res1[3255],mul_res1[3256],mul_res1[3257],mul_res1[3258],mul_res1[3259],mul_res1[3260],mul_res1[3261],mul_res1[3262],mul_res1[3263],mul_res1[3264],mul_res1[3265],mul_res1[3266],mul_res1[3267],mul_res1[3268],mul_res1[3269],mul_res1[3270],mul_res1[3271],mul_res1[3272],mul_res1[3273],mul_res1[3274],mul_res1[3275],mul_res1[3276],mul_res1[3277],mul_res1[3278],mul_res1[3279],mul_res1[3280],mul_res1[3281],mul_res1[3282],mul_res1[3283],mul_res1[3284],mul_res1[3285],mul_res1[3286],mul_res1[3287],mul_res1[3288],mul_res1[3289],mul_res1[3290],mul_res1[3291],mul_res1[3292],mul_res1[3293],mul_res1[3294],mul_res1[3295],mul_res1[3296],mul_res1[3297],mul_res1[3298],mul_res1[3299],mul_res1[3300],mul_res1[3301],mul_res1[3302],mul_res1[3303],mul_res1[3304],mul_res1[3305],mul_res1[3306],mul_res1[3307],mul_res1[3308],mul_res1[3309],mul_res1[3310],mul_res1[3311],mul_res1[3312],mul_res1[3313],mul_res1[3314],mul_res1[3315],mul_res1[3316],mul_res1[3317],mul_res1[3318],mul_res1[3319],mul_res1[3320],mul_res1[3321],mul_res1[3322],mul_res1[3323],mul_res1[3324],mul_res1[3325],mul_res1[3326],mul_res1[3327],mul_res1[3328],mul_res1[3329],mul_res1[3330],mul_res1[3331],mul_res1[3332],mul_res1[3333],mul_res1[3334],mul_res1[3335],mul_res1[3336],mul_res1[3337],mul_res1[3338],mul_res1[3339],mul_res1[3340],mul_res1[3341],mul_res1[3342],mul_res1[3343],mul_res1[3344],mul_res1[3345],mul_res1[3346],mul_res1[3347],mul_res1[3348],mul_res1[3349],mul_res1[3350],mul_res1[3351],mul_res1[3352],mul_res1[3353],mul_res1[3354],mul_res1[3355],mul_res1[3356],mul_res1[3357],mul_res1[3358],mul_res1[3359],mul_res1[3360],mul_res1[3361],mul_res1[3362],mul_res1[3363],mul_res1[3364],mul_res1[3365],mul_res1[3366],mul_res1[3367],mul_res1[3368],mul_res1[3369],mul_res1[3370],mul_res1[3371],mul_res1[3372],mul_res1[3373],mul_res1[3374],mul_res1[3375],mul_res1[3376],mul_res1[3377],mul_res1[3378],mul_res1[3379],mul_res1[3380],mul_res1[3381],mul_res1[3382],mul_res1[3383],mul_res1[3384],mul_res1[3385],mul_res1[3386],mul_res1[3387],mul_res1[3388],mul_res1[3389],mul_res1[3390],mul_res1[3391],mul_res1[3392],mul_res1[3393],mul_res1[3394],mul_res1[3395],mul_res1[3396],mul_res1[3397],mul_res1[3398],mul_res1[3399],result_fc1[16]);


adder_200in adder_200in_mod_17(clk,rst,mul_res1[3400],mul_res1[3401],mul_res1[3402],mul_res1[3403],mul_res1[3404],mul_res1[3405],mul_res1[3406],mul_res1[3407],mul_res1[3408],mul_res1[3409],mul_res1[3410],mul_res1[3411],mul_res1[3412],mul_res1[3413],mul_res1[3414],mul_res1[3415],mul_res1[3416],mul_res1[3417],mul_res1[3418],mul_res1[3419],mul_res1[3420],mul_res1[3421],mul_res1[3422],mul_res1[3423],mul_res1[3424],mul_res1[3425],mul_res1[3426],mul_res1[3427],mul_res1[3428],mul_res1[3429],mul_res1[3430],mul_res1[3431],mul_res1[3432],mul_res1[3433],mul_res1[3434],mul_res1[3435],mul_res1[3436],mul_res1[3437],mul_res1[3438],mul_res1[3439],mul_res1[3440],mul_res1[3441],mul_res1[3442],mul_res1[3443],mul_res1[3444],mul_res1[3445],mul_res1[3446],mul_res1[3447],mul_res1[3448],mul_res1[3449],mul_res1[3450],mul_res1[3451],mul_res1[3452],mul_res1[3453],mul_res1[3454],mul_res1[3455],mul_res1[3456],mul_res1[3457],mul_res1[3458],mul_res1[3459],mul_res1[3460],mul_res1[3461],mul_res1[3462],mul_res1[3463],mul_res1[3464],mul_res1[3465],mul_res1[3466],mul_res1[3467],mul_res1[3468],mul_res1[3469],mul_res1[3470],mul_res1[3471],mul_res1[3472],mul_res1[3473],mul_res1[3474],mul_res1[3475],mul_res1[3476],mul_res1[3477],mul_res1[3478],mul_res1[3479],mul_res1[3480],mul_res1[3481],mul_res1[3482],mul_res1[3483],mul_res1[3484],mul_res1[3485],mul_res1[3486],mul_res1[3487],mul_res1[3488],mul_res1[3489],mul_res1[3490],mul_res1[3491],mul_res1[3492],mul_res1[3493],mul_res1[3494],mul_res1[3495],mul_res1[3496],mul_res1[3497],mul_res1[3498],mul_res1[3499],mul_res1[3500],mul_res1[3501],mul_res1[3502],mul_res1[3503],mul_res1[3504],mul_res1[3505],mul_res1[3506],mul_res1[3507],mul_res1[3508],mul_res1[3509],mul_res1[3510],mul_res1[3511],mul_res1[3512],mul_res1[3513],mul_res1[3514],mul_res1[3515],mul_res1[3516],mul_res1[3517],mul_res1[3518],mul_res1[3519],mul_res1[3520],mul_res1[3521],mul_res1[3522],mul_res1[3523],mul_res1[3524],mul_res1[3525],mul_res1[3526],mul_res1[3527],mul_res1[3528],mul_res1[3529],mul_res1[3530],mul_res1[3531],mul_res1[3532],mul_res1[3533],mul_res1[3534],mul_res1[3535],mul_res1[3536],mul_res1[3537],mul_res1[3538],mul_res1[3539],mul_res1[3540],mul_res1[3541],mul_res1[3542],mul_res1[3543],mul_res1[3544],mul_res1[3545],mul_res1[3546],mul_res1[3547],mul_res1[3548],mul_res1[3549],mul_res1[3550],mul_res1[3551],mul_res1[3552],mul_res1[3553],mul_res1[3554],mul_res1[3555],mul_res1[3556],mul_res1[3557],mul_res1[3558],mul_res1[3559],mul_res1[3560],mul_res1[3561],mul_res1[3562],mul_res1[3563],mul_res1[3564],mul_res1[3565],mul_res1[3566],mul_res1[3567],mul_res1[3568],mul_res1[3569],mul_res1[3570],mul_res1[3571],mul_res1[3572],mul_res1[3573],mul_res1[3574],mul_res1[3575],mul_res1[3576],mul_res1[3577],mul_res1[3578],mul_res1[3579],mul_res1[3580],mul_res1[3581],mul_res1[3582],mul_res1[3583],mul_res1[3584],mul_res1[3585],mul_res1[3586],mul_res1[3587],mul_res1[3588],mul_res1[3589],mul_res1[3590],mul_res1[3591],mul_res1[3592],mul_res1[3593],mul_res1[3594],mul_res1[3595],mul_res1[3596],mul_res1[3597],mul_res1[3598],mul_res1[3599],result_fc1[17]);


adder_200in adder_200in_mod_18(clk,rst,mul_res1[3600],mul_res1[3601],mul_res1[3602],mul_res1[3603],mul_res1[3604],mul_res1[3605],mul_res1[3606],mul_res1[3607],mul_res1[3608],mul_res1[3609],mul_res1[3610],mul_res1[3611],mul_res1[3612],mul_res1[3613],mul_res1[3614],mul_res1[3615],mul_res1[3616],mul_res1[3617],mul_res1[3618],mul_res1[3619],mul_res1[3620],mul_res1[3621],mul_res1[3622],mul_res1[3623],mul_res1[3624],mul_res1[3625],mul_res1[3626],mul_res1[3627],mul_res1[3628],mul_res1[3629],mul_res1[3630],mul_res1[3631],mul_res1[3632],mul_res1[3633],mul_res1[3634],mul_res1[3635],mul_res1[3636],mul_res1[3637],mul_res1[3638],mul_res1[3639],mul_res1[3640],mul_res1[3641],mul_res1[3642],mul_res1[3643],mul_res1[3644],mul_res1[3645],mul_res1[3646],mul_res1[3647],mul_res1[3648],mul_res1[3649],mul_res1[3650],mul_res1[3651],mul_res1[3652],mul_res1[3653],mul_res1[3654],mul_res1[3655],mul_res1[3656],mul_res1[3657],mul_res1[3658],mul_res1[3659],mul_res1[3660],mul_res1[3661],mul_res1[3662],mul_res1[3663],mul_res1[3664],mul_res1[3665],mul_res1[3666],mul_res1[3667],mul_res1[3668],mul_res1[3669],mul_res1[3670],mul_res1[3671],mul_res1[3672],mul_res1[3673],mul_res1[3674],mul_res1[3675],mul_res1[3676],mul_res1[3677],mul_res1[3678],mul_res1[3679],mul_res1[3680],mul_res1[3681],mul_res1[3682],mul_res1[3683],mul_res1[3684],mul_res1[3685],mul_res1[3686],mul_res1[3687],mul_res1[3688],mul_res1[3689],mul_res1[3690],mul_res1[3691],mul_res1[3692],mul_res1[3693],mul_res1[3694],mul_res1[3695],mul_res1[3696],mul_res1[3697],mul_res1[3698],mul_res1[3699],mul_res1[3700],mul_res1[3701],mul_res1[3702],mul_res1[3703],mul_res1[3704],mul_res1[3705],mul_res1[3706],mul_res1[3707],mul_res1[3708],mul_res1[3709],mul_res1[3710],mul_res1[3711],mul_res1[3712],mul_res1[3713],mul_res1[3714],mul_res1[3715],mul_res1[3716],mul_res1[3717],mul_res1[3718],mul_res1[3719],mul_res1[3720],mul_res1[3721],mul_res1[3722],mul_res1[3723],mul_res1[3724],mul_res1[3725],mul_res1[3726],mul_res1[3727],mul_res1[3728],mul_res1[3729],mul_res1[3730],mul_res1[3731],mul_res1[3732],mul_res1[3733],mul_res1[3734],mul_res1[3735],mul_res1[3736],mul_res1[3737],mul_res1[3738],mul_res1[3739],mul_res1[3740],mul_res1[3741],mul_res1[3742],mul_res1[3743],mul_res1[3744],mul_res1[3745],mul_res1[3746],mul_res1[3747],mul_res1[3748],mul_res1[3749],mul_res1[3750],mul_res1[3751],mul_res1[3752],mul_res1[3753],mul_res1[3754],mul_res1[3755],mul_res1[3756],mul_res1[3757],mul_res1[3758],mul_res1[3759],mul_res1[3760],mul_res1[3761],mul_res1[3762],mul_res1[3763],mul_res1[3764],mul_res1[3765],mul_res1[3766],mul_res1[3767],mul_res1[3768],mul_res1[3769],mul_res1[3770],mul_res1[3771],mul_res1[3772],mul_res1[3773],mul_res1[3774],mul_res1[3775],mul_res1[3776],mul_res1[3777],mul_res1[3778],mul_res1[3779],mul_res1[3780],mul_res1[3781],mul_res1[3782],mul_res1[3783],mul_res1[3784],mul_res1[3785],mul_res1[3786],mul_res1[3787],mul_res1[3788],mul_res1[3789],mul_res1[3790],mul_res1[3791],mul_res1[3792],mul_res1[3793],mul_res1[3794],mul_res1[3795],mul_res1[3796],mul_res1[3797],mul_res1[3798],mul_res1[3799],result_fc1[18]);


adder_200in adder_200in_mod_19(clk,rst,mul_res1[3800],mul_res1[3801],mul_res1[3802],mul_res1[3803],mul_res1[3804],mul_res1[3805],mul_res1[3806],mul_res1[3807],mul_res1[3808],mul_res1[3809],mul_res1[3810],mul_res1[3811],mul_res1[3812],mul_res1[3813],mul_res1[3814],mul_res1[3815],mul_res1[3816],mul_res1[3817],mul_res1[3818],mul_res1[3819],mul_res1[3820],mul_res1[3821],mul_res1[3822],mul_res1[3823],mul_res1[3824],mul_res1[3825],mul_res1[3826],mul_res1[3827],mul_res1[3828],mul_res1[3829],mul_res1[3830],mul_res1[3831],mul_res1[3832],mul_res1[3833],mul_res1[3834],mul_res1[3835],mul_res1[3836],mul_res1[3837],mul_res1[3838],mul_res1[3839],mul_res1[3840],mul_res1[3841],mul_res1[3842],mul_res1[3843],mul_res1[3844],mul_res1[3845],mul_res1[3846],mul_res1[3847],mul_res1[3848],mul_res1[3849],mul_res1[3850],mul_res1[3851],mul_res1[3852],mul_res1[3853],mul_res1[3854],mul_res1[3855],mul_res1[3856],mul_res1[3857],mul_res1[3858],mul_res1[3859],mul_res1[3860],mul_res1[3861],mul_res1[3862],mul_res1[3863],mul_res1[3864],mul_res1[3865],mul_res1[3866],mul_res1[3867],mul_res1[3868],mul_res1[3869],mul_res1[3870],mul_res1[3871],mul_res1[3872],mul_res1[3873],mul_res1[3874],mul_res1[3875],mul_res1[3876],mul_res1[3877],mul_res1[3878],mul_res1[3879],mul_res1[3880],mul_res1[3881],mul_res1[3882],mul_res1[3883],mul_res1[3884],mul_res1[3885],mul_res1[3886],mul_res1[3887],mul_res1[3888],mul_res1[3889],mul_res1[3890],mul_res1[3891],mul_res1[3892],mul_res1[3893],mul_res1[3894],mul_res1[3895],mul_res1[3896],mul_res1[3897],mul_res1[3898],mul_res1[3899],mul_res1[3900],mul_res1[3901],mul_res1[3902],mul_res1[3903],mul_res1[3904],mul_res1[3905],mul_res1[3906],mul_res1[3907],mul_res1[3908],mul_res1[3909],mul_res1[3910],mul_res1[3911],mul_res1[3912],mul_res1[3913],mul_res1[3914],mul_res1[3915],mul_res1[3916],mul_res1[3917],mul_res1[3918],mul_res1[3919],mul_res1[3920],mul_res1[3921],mul_res1[3922],mul_res1[3923],mul_res1[3924],mul_res1[3925],mul_res1[3926],mul_res1[3927],mul_res1[3928],mul_res1[3929],mul_res1[3930],mul_res1[3931],mul_res1[3932],mul_res1[3933],mul_res1[3934],mul_res1[3935],mul_res1[3936],mul_res1[3937],mul_res1[3938],mul_res1[3939],mul_res1[3940],mul_res1[3941],mul_res1[3942],mul_res1[3943],mul_res1[3944],mul_res1[3945],mul_res1[3946],mul_res1[3947],mul_res1[3948],mul_res1[3949],mul_res1[3950],mul_res1[3951],mul_res1[3952],mul_res1[3953],mul_res1[3954],mul_res1[3955],mul_res1[3956],mul_res1[3957],mul_res1[3958],mul_res1[3959],mul_res1[3960],mul_res1[3961],mul_res1[3962],mul_res1[3963],mul_res1[3964],mul_res1[3965],mul_res1[3966],mul_res1[3967],mul_res1[3968],mul_res1[3969],mul_res1[3970],mul_res1[3971],mul_res1[3972],mul_res1[3973],mul_res1[3974],mul_res1[3975],mul_res1[3976],mul_res1[3977],mul_res1[3978],mul_res1[3979],mul_res1[3980],mul_res1[3981],mul_res1[3982],mul_res1[3983],mul_res1[3984],mul_res1[3985],mul_res1[3986],mul_res1[3987],mul_res1[3988],mul_res1[3989],mul_res1[3990],mul_res1[3991],mul_res1[3992],mul_res1[3993],mul_res1[3994],mul_res1[3995],mul_res1[3996],mul_res1[3997],mul_res1[3998],mul_res1[3999],result_fc1[19]);


adder_200in adder_200in_mod_20(clk,rst,mul_res1[4000],mul_res1[4001],mul_res1[4002],mul_res1[4003],mul_res1[4004],mul_res1[4005],mul_res1[4006],mul_res1[4007],mul_res1[4008],mul_res1[4009],mul_res1[4010],mul_res1[4011],mul_res1[4012],mul_res1[4013],mul_res1[4014],mul_res1[4015],mul_res1[4016],mul_res1[4017],mul_res1[4018],mul_res1[4019],mul_res1[4020],mul_res1[4021],mul_res1[4022],mul_res1[4023],mul_res1[4024],mul_res1[4025],mul_res1[4026],mul_res1[4027],mul_res1[4028],mul_res1[4029],mul_res1[4030],mul_res1[4031],mul_res1[4032],mul_res1[4033],mul_res1[4034],mul_res1[4035],mul_res1[4036],mul_res1[4037],mul_res1[4038],mul_res1[4039],mul_res1[4040],mul_res1[4041],mul_res1[4042],mul_res1[4043],mul_res1[4044],mul_res1[4045],mul_res1[4046],mul_res1[4047],mul_res1[4048],mul_res1[4049],mul_res1[4050],mul_res1[4051],mul_res1[4052],mul_res1[4053],mul_res1[4054],mul_res1[4055],mul_res1[4056],mul_res1[4057],mul_res1[4058],mul_res1[4059],mul_res1[4060],mul_res1[4061],mul_res1[4062],mul_res1[4063],mul_res1[4064],mul_res1[4065],mul_res1[4066],mul_res1[4067],mul_res1[4068],mul_res1[4069],mul_res1[4070],mul_res1[4071],mul_res1[4072],mul_res1[4073],mul_res1[4074],mul_res1[4075],mul_res1[4076],mul_res1[4077],mul_res1[4078],mul_res1[4079],mul_res1[4080],mul_res1[4081],mul_res1[4082],mul_res1[4083],mul_res1[4084],mul_res1[4085],mul_res1[4086],mul_res1[4087],mul_res1[4088],mul_res1[4089],mul_res1[4090],mul_res1[4091],mul_res1[4092],mul_res1[4093],mul_res1[4094],mul_res1[4095],mul_res1[4096],mul_res1[4097],mul_res1[4098],mul_res1[4099],mul_res1[4100],mul_res1[4101],mul_res1[4102],mul_res1[4103],mul_res1[4104],mul_res1[4105],mul_res1[4106],mul_res1[4107],mul_res1[4108],mul_res1[4109],mul_res1[4110],mul_res1[4111],mul_res1[4112],mul_res1[4113],mul_res1[4114],mul_res1[4115],mul_res1[4116],mul_res1[4117],mul_res1[4118],mul_res1[4119],mul_res1[4120],mul_res1[4121],mul_res1[4122],mul_res1[4123],mul_res1[4124],mul_res1[4125],mul_res1[4126],mul_res1[4127],mul_res1[4128],mul_res1[4129],mul_res1[4130],mul_res1[4131],mul_res1[4132],mul_res1[4133],mul_res1[4134],mul_res1[4135],mul_res1[4136],mul_res1[4137],mul_res1[4138],mul_res1[4139],mul_res1[4140],mul_res1[4141],mul_res1[4142],mul_res1[4143],mul_res1[4144],mul_res1[4145],mul_res1[4146],mul_res1[4147],mul_res1[4148],mul_res1[4149],mul_res1[4150],mul_res1[4151],mul_res1[4152],mul_res1[4153],mul_res1[4154],mul_res1[4155],mul_res1[4156],mul_res1[4157],mul_res1[4158],mul_res1[4159],mul_res1[4160],mul_res1[4161],mul_res1[4162],mul_res1[4163],mul_res1[4164],mul_res1[4165],mul_res1[4166],mul_res1[4167],mul_res1[4168],mul_res1[4169],mul_res1[4170],mul_res1[4171],mul_res1[4172],mul_res1[4173],mul_res1[4174],mul_res1[4175],mul_res1[4176],mul_res1[4177],mul_res1[4178],mul_res1[4179],mul_res1[4180],mul_res1[4181],mul_res1[4182],mul_res1[4183],mul_res1[4184],mul_res1[4185],mul_res1[4186],mul_res1[4187],mul_res1[4188],mul_res1[4189],mul_res1[4190],mul_res1[4191],mul_res1[4192],mul_res1[4193],mul_res1[4194],mul_res1[4195],mul_res1[4196],mul_res1[4197],mul_res1[4198],mul_res1[4199],result_fc1[20]);


adder_200in adder_200in_mod_21(clk,rst,mul_res1[4200],mul_res1[4201],mul_res1[4202],mul_res1[4203],mul_res1[4204],mul_res1[4205],mul_res1[4206],mul_res1[4207],mul_res1[4208],mul_res1[4209],mul_res1[4210],mul_res1[4211],mul_res1[4212],mul_res1[4213],mul_res1[4214],mul_res1[4215],mul_res1[4216],mul_res1[4217],mul_res1[4218],mul_res1[4219],mul_res1[4220],mul_res1[4221],mul_res1[4222],mul_res1[4223],mul_res1[4224],mul_res1[4225],mul_res1[4226],mul_res1[4227],mul_res1[4228],mul_res1[4229],mul_res1[4230],mul_res1[4231],mul_res1[4232],mul_res1[4233],mul_res1[4234],mul_res1[4235],mul_res1[4236],mul_res1[4237],mul_res1[4238],mul_res1[4239],mul_res1[4240],mul_res1[4241],mul_res1[4242],mul_res1[4243],mul_res1[4244],mul_res1[4245],mul_res1[4246],mul_res1[4247],mul_res1[4248],mul_res1[4249],mul_res1[4250],mul_res1[4251],mul_res1[4252],mul_res1[4253],mul_res1[4254],mul_res1[4255],mul_res1[4256],mul_res1[4257],mul_res1[4258],mul_res1[4259],mul_res1[4260],mul_res1[4261],mul_res1[4262],mul_res1[4263],mul_res1[4264],mul_res1[4265],mul_res1[4266],mul_res1[4267],mul_res1[4268],mul_res1[4269],mul_res1[4270],mul_res1[4271],mul_res1[4272],mul_res1[4273],mul_res1[4274],mul_res1[4275],mul_res1[4276],mul_res1[4277],mul_res1[4278],mul_res1[4279],mul_res1[4280],mul_res1[4281],mul_res1[4282],mul_res1[4283],mul_res1[4284],mul_res1[4285],mul_res1[4286],mul_res1[4287],mul_res1[4288],mul_res1[4289],mul_res1[4290],mul_res1[4291],mul_res1[4292],mul_res1[4293],mul_res1[4294],mul_res1[4295],mul_res1[4296],mul_res1[4297],mul_res1[4298],mul_res1[4299],mul_res1[4300],mul_res1[4301],mul_res1[4302],mul_res1[4303],mul_res1[4304],mul_res1[4305],mul_res1[4306],mul_res1[4307],mul_res1[4308],mul_res1[4309],mul_res1[4310],mul_res1[4311],mul_res1[4312],mul_res1[4313],mul_res1[4314],mul_res1[4315],mul_res1[4316],mul_res1[4317],mul_res1[4318],mul_res1[4319],mul_res1[4320],mul_res1[4321],mul_res1[4322],mul_res1[4323],mul_res1[4324],mul_res1[4325],mul_res1[4326],mul_res1[4327],mul_res1[4328],mul_res1[4329],mul_res1[4330],mul_res1[4331],mul_res1[4332],mul_res1[4333],mul_res1[4334],mul_res1[4335],mul_res1[4336],mul_res1[4337],mul_res1[4338],mul_res1[4339],mul_res1[4340],mul_res1[4341],mul_res1[4342],mul_res1[4343],mul_res1[4344],mul_res1[4345],mul_res1[4346],mul_res1[4347],mul_res1[4348],mul_res1[4349],mul_res1[4350],mul_res1[4351],mul_res1[4352],mul_res1[4353],mul_res1[4354],mul_res1[4355],mul_res1[4356],mul_res1[4357],mul_res1[4358],mul_res1[4359],mul_res1[4360],mul_res1[4361],mul_res1[4362],mul_res1[4363],mul_res1[4364],mul_res1[4365],mul_res1[4366],mul_res1[4367],mul_res1[4368],mul_res1[4369],mul_res1[4370],mul_res1[4371],mul_res1[4372],mul_res1[4373],mul_res1[4374],mul_res1[4375],mul_res1[4376],mul_res1[4377],mul_res1[4378],mul_res1[4379],mul_res1[4380],mul_res1[4381],mul_res1[4382],mul_res1[4383],mul_res1[4384],mul_res1[4385],mul_res1[4386],mul_res1[4387],mul_res1[4388],mul_res1[4389],mul_res1[4390],mul_res1[4391],mul_res1[4392],mul_res1[4393],mul_res1[4394],mul_res1[4395],mul_res1[4396],mul_res1[4397],mul_res1[4398],mul_res1[4399],result_fc1[21]);


adder_200in adder_200in_mod_22(clk,rst,mul_res1[4400],mul_res1[4401],mul_res1[4402],mul_res1[4403],mul_res1[4404],mul_res1[4405],mul_res1[4406],mul_res1[4407],mul_res1[4408],mul_res1[4409],mul_res1[4410],mul_res1[4411],mul_res1[4412],mul_res1[4413],mul_res1[4414],mul_res1[4415],mul_res1[4416],mul_res1[4417],mul_res1[4418],mul_res1[4419],mul_res1[4420],mul_res1[4421],mul_res1[4422],mul_res1[4423],mul_res1[4424],mul_res1[4425],mul_res1[4426],mul_res1[4427],mul_res1[4428],mul_res1[4429],mul_res1[4430],mul_res1[4431],mul_res1[4432],mul_res1[4433],mul_res1[4434],mul_res1[4435],mul_res1[4436],mul_res1[4437],mul_res1[4438],mul_res1[4439],mul_res1[4440],mul_res1[4441],mul_res1[4442],mul_res1[4443],mul_res1[4444],mul_res1[4445],mul_res1[4446],mul_res1[4447],mul_res1[4448],mul_res1[4449],mul_res1[4450],mul_res1[4451],mul_res1[4452],mul_res1[4453],mul_res1[4454],mul_res1[4455],mul_res1[4456],mul_res1[4457],mul_res1[4458],mul_res1[4459],mul_res1[4460],mul_res1[4461],mul_res1[4462],mul_res1[4463],mul_res1[4464],mul_res1[4465],mul_res1[4466],mul_res1[4467],mul_res1[4468],mul_res1[4469],mul_res1[4470],mul_res1[4471],mul_res1[4472],mul_res1[4473],mul_res1[4474],mul_res1[4475],mul_res1[4476],mul_res1[4477],mul_res1[4478],mul_res1[4479],mul_res1[4480],mul_res1[4481],mul_res1[4482],mul_res1[4483],mul_res1[4484],mul_res1[4485],mul_res1[4486],mul_res1[4487],mul_res1[4488],mul_res1[4489],mul_res1[4490],mul_res1[4491],mul_res1[4492],mul_res1[4493],mul_res1[4494],mul_res1[4495],mul_res1[4496],mul_res1[4497],mul_res1[4498],mul_res1[4499],mul_res1[4500],mul_res1[4501],mul_res1[4502],mul_res1[4503],mul_res1[4504],mul_res1[4505],mul_res1[4506],mul_res1[4507],mul_res1[4508],mul_res1[4509],mul_res1[4510],mul_res1[4511],mul_res1[4512],mul_res1[4513],mul_res1[4514],mul_res1[4515],mul_res1[4516],mul_res1[4517],mul_res1[4518],mul_res1[4519],mul_res1[4520],mul_res1[4521],mul_res1[4522],mul_res1[4523],mul_res1[4524],mul_res1[4525],mul_res1[4526],mul_res1[4527],mul_res1[4528],mul_res1[4529],mul_res1[4530],mul_res1[4531],mul_res1[4532],mul_res1[4533],mul_res1[4534],mul_res1[4535],mul_res1[4536],mul_res1[4537],mul_res1[4538],mul_res1[4539],mul_res1[4540],mul_res1[4541],mul_res1[4542],mul_res1[4543],mul_res1[4544],mul_res1[4545],mul_res1[4546],mul_res1[4547],mul_res1[4548],mul_res1[4549],mul_res1[4550],mul_res1[4551],mul_res1[4552],mul_res1[4553],mul_res1[4554],mul_res1[4555],mul_res1[4556],mul_res1[4557],mul_res1[4558],mul_res1[4559],mul_res1[4560],mul_res1[4561],mul_res1[4562],mul_res1[4563],mul_res1[4564],mul_res1[4565],mul_res1[4566],mul_res1[4567],mul_res1[4568],mul_res1[4569],mul_res1[4570],mul_res1[4571],mul_res1[4572],mul_res1[4573],mul_res1[4574],mul_res1[4575],mul_res1[4576],mul_res1[4577],mul_res1[4578],mul_res1[4579],mul_res1[4580],mul_res1[4581],mul_res1[4582],mul_res1[4583],mul_res1[4584],mul_res1[4585],mul_res1[4586],mul_res1[4587],mul_res1[4588],mul_res1[4589],mul_res1[4590],mul_res1[4591],mul_res1[4592],mul_res1[4593],mul_res1[4594],mul_res1[4595],mul_res1[4596],mul_res1[4597],mul_res1[4598],mul_res1[4599],result_fc1[22]);


adder_200in adder_200in_mod_23(clk,rst,mul_res1[4600],mul_res1[4601],mul_res1[4602],mul_res1[4603],mul_res1[4604],mul_res1[4605],mul_res1[4606],mul_res1[4607],mul_res1[4608],mul_res1[4609],mul_res1[4610],mul_res1[4611],mul_res1[4612],mul_res1[4613],mul_res1[4614],mul_res1[4615],mul_res1[4616],mul_res1[4617],mul_res1[4618],mul_res1[4619],mul_res1[4620],mul_res1[4621],mul_res1[4622],mul_res1[4623],mul_res1[4624],mul_res1[4625],mul_res1[4626],mul_res1[4627],mul_res1[4628],mul_res1[4629],mul_res1[4630],mul_res1[4631],mul_res1[4632],mul_res1[4633],mul_res1[4634],mul_res1[4635],mul_res1[4636],mul_res1[4637],mul_res1[4638],mul_res1[4639],mul_res1[4640],mul_res1[4641],mul_res1[4642],mul_res1[4643],mul_res1[4644],mul_res1[4645],mul_res1[4646],mul_res1[4647],mul_res1[4648],mul_res1[4649],mul_res1[4650],mul_res1[4651],mul_res1[4652],mul_res1[4653],mul_res1[4654],mul_res1[4655],mul_res1[4656],mul_res1[4657],mul_res1[4658],mul_res1[4659],mul_res1[4660],mul_res1[4661],mul_res1[4662],mul_res1[4663],mul_res1[4664],mul_res1[4665],mul_res1[4666],mul_res1[4667],mul_res1[4668],mul_res1[4669],mul_res1[4670],mul_res1[4671],mul_res1[4672],mul_res1[4673],mul_res1[4674],mul_res1[4675],mul_res1[4676],mul_res1[4677],mul_res1[4678],mul_res1[4679],mul_res1[4680],mul_res1[4681],mul_res1[4682],mul_res1[4683],mul_res1[4684],mul_res1[4685],mul_res1[4686],mul_res1[4687],mul_res1[4688],mul_res1[4689],mul_res1[4690],mul_res1[4691],mul_res1[4692],mul_res1[4693],mul_res1[4694],mul_res1[4695],mul_res1[4696],mul_res1[4697],mul_res1[4698],mul_res1[4699],mul_res1[4700],mul_res1[4701],mul_res1[4702],mul_res1[4703],mul_res1[4704],mul_res1[4705],mul_res1[4706],mul_res1[4707],mul_res1[4708],mul_res1[4709],mul_res1[4710],mul_res1[4711],mul_res1[4712],mul_res1[4713],mul_res1[4714],mul_res1[4715],mul_res1[4716],mul_res1[4717],mul_res1[4718],mul_res1[4719],mul_res1[4720],mul_res1[4721],mul_res1[4722],mul_res1[4723],mul_res1[4724],mul_res1[4725],mul_res1[4726],mul_res1[4727],mul_res1[4728],mul_res1[4729],mul_res1[4730],mul_res1[4731],mul_res1[4732],mul_res1[4733],mul_res1[4734],mul_res1[4735],mul_res1[4736],mul_res1[4737],mul_res1[4738],mul_res1[4739],mul_res1[4740],mul_res1[4741],mul_res1[4742],mul_res1[4743],mul_res1[4744],mul_res1[4745],mul_res1[4746],mul_res1[4747],mul_res1[4748],mul_res1[4749],mul_res1[4750],mul_res1[4751],mul_res1[4752],mul_res1[4753],mul_res1[4754],mul_res1[4755],mul_res1[4756],mul_res1[4757],mul_res1[4758],mul_res1[4759],mul_res1[4760],mul_res1[4761],mul_res1[4762],mul_res1[4763],mul_res1[4764],mul_res1[4765],mul_res1[4766],mul_res1[4767],mul_res1[4768],mul_res1[4769],mul_res1[4770],mul_res1[4771],mul_res1[4772],mul_res1[4773],mul_res1[4774],mul_res1[4775],mul_res1[4776],mul_res1[4777],mul_res1[4778],mul_res1[4779],mul_res1[4780],mul_res1[4781],mul_res1[4782],mul_res1[4783],mul_res1[4784],mul_res1[4785],mul_res1[4786],mul_res1[4787],mul_res1[4788],mul_res1[4789],mul_res1[4790],mul_res1[4791],mul_res1[4792],mul_res1[4793],mul_res1[4794],mul_res1[4795],mul_res1[4796],mul_res1[4797],mul_res1[4798],mul_res1[4799],result_fc1[23]);


adder_200in adder_200in_mod_24(clk,rst,mul_res1[4800],mul_res1[4801],mul_res1[4802],mul_res1[4803],mul_res1[4804],mul_res1[4805],mul_res1[4806],mul_res1[4807],mul_res1[4808],mul_res1[4809],mul_res1[4810],mul_res1[4811],mul_res1[4812],mul_res1[4813],mul_res1[4814],mul_res1[4815],mul_res1[4816],mul_res1[4817],mul_res1[4818],mul_res1[4819],mul_res1[4820],mul_res1[4821],mul_res1[4822],mul_res1[4823],mul_res1[4824],mul_res1[4825],mul_res1[4826],mul_res1[4827],mul_res1[4828],mul_res1[4829],mul_res1[4830],mul_res1[4831],mul_res1[4832],mul_res1[4833],mul_res1[4834],mul_res1[4835],mul_res1[4836],mul_res1[4837],mul_res1[4838],mul_res1[4839],mul_res1[4840],mul_res1[4841],mul_res1[4842],mul_res1[4843],mul_res1[4844],mul_res1[4845],mul_res1[4846],mul_res1[4847],mul_res1[4848],mul_res1[4849],mul_res1[4850],mul_res1[4851],mul_res1[4852],mul_res1[4853],mul_res1[4854],mul_res1[4855],mul_res1[4856],mul_res1[4857],mul_res1[4858],mul_res1[4859],mul_res1[4860],mul_res1[4861],mul_res1[4862],mul_res1[4863],mul_res1[4864],mul_res1[4865],mul_res1[4866],mul_res1[4867],mul_res1[4868],mul_res1[4869],mul_res1[4870],mul_res1[4871],mul_res1[4872],mul_res1[4873],mul_res1[4874],mul_res1[4875],mul_res1[4876],mul_res1[4877],mul_res1[4878],mul_res1[4879],mul_res1[4880],mul_res1[4881],mul_res1[4882],mul_res1[4883],mul_res1[4884],mul_res1[4885],mul_res1[4886],mul_res1[4887],mul_res1[4888],mul_res1[4889],mul_res1[4890],mul_res1[4891],mul_res1[4892],mul_res1[4893],mul_res1[4894],mul_res1[4895],mul_res1[4896],mul_res1[4897],mul_res1[4898],mul_res1[4899],mul_res1[4900],mul_res1[4901],mul_res1[4902],mul_res1[4903],mul_res1[4904],mul_res1[4905],mul_res1[4906],mul_res1[4907],mul_res1[4908],mul_res1[4909],mul_res1[4910],mul_res1[4911],mul_res1[4912],mul_res1[4913],mul_res1[4914],mul_res1[4915],mul_res1[4916],mul_res1[4917],mul_res1[4918],mul_res1[4919],mul_res1[4920],mul_res1[4921],mul_res1[4922],mul_res1[4923],mul_res1[4924],mul_res1[4925],mul_res1[4926],mul_res1[4927],mul_res1[4928],mul_res1[4929],mul_res1[4930],mul_res1[4931],mul_res1[4932],mul_res1[4933],mul_res1[4934],mul_res1[4935],mul_res1[4936],mul_res1[4937],mul_res1[4938],mul_res1[4939],mul_res1[4940],mul_res1[4941],mul_res1[4942],mul_res1[4943],mul_res1[4944],mul_res1[4945],mul_res1[4946],mul_res1[4947],mul_res1[4948],mul_res1[4949],mul_res1[4950],mul_res1[4951],mul_res1[4952],mul_res1[4953],mul_res1[4954],mul_res1[4955],mul_res1[4956],mul_res1[4957],mul_res1[4958],mul_res1[4959],mul_res1[4960],mul_res1[4961],mul_res1[4962],mul_res1[4963],mul_res1[4964],mul_res1[4965],mul_res1[4966],mul_res1[4967],mul_res1[4968],mul_res1[4969],mul_res1[4970],mul_res1[4971],mul_res1[4972],mul_res1[4973],mul_res1[4974],mul_res1[4975],mul_res1[4976],mul_res1[4977],mul_res1[4978],mul_res1[4979],mul_res1[4980],mul_res1[4981],mul_res1[4982],mul_res1[4983],mul_res1[4984],mul_res1[4985],mul_res1[4986],mul_res1[4987],mul_res1[4988],mul_res1[4989],mul_res1[4990],mul_res1[4991],mul_res1[4992],mul_res1[4993],mul_res1[4994],mul_res1[4995],mul_res1[4996],mul_res1[4997],mul_res1[4998],mul_res1[4999],result_fc1[24]);


adder_200in adder_200in_mod_25(clk,rst,mul_res1[5000],mul_res1[5001],mul_res1[5002],mul_res1[5003],mul_res1[5004],mul_res1[5005],mul_res1[5006],mul_res1[5007],mul_res1[5008],mul_res1[5009],mul_res1[5010],mul_res1[5011],mul_res1[5012],mul_res1[5013],mul_res1[5014],mul_res1[5015],mul_res1[5016],mul_res1[5017],mul_res1[5018],mul_res1[5019],mul_res1[5020],mul_res1[5021],mul_res1[5022],mul_res1[5023],mul_res1[5024],mul_res1[5025],mul_res1[5026],mul_res1[5027],mul_res1[5028],mul_res1[5029],mul_res1[5030],mul_res1[5031],mul_res1[5032],mul_res1[5033],mul_res1[5034],mul_res1[5035],mul_res1[5036],mul_res1[5037],mul_res1[5038],mul_res1[5039],mul_res1[5040],mul_res1[5041],mul_res1[5042],mul_res1[5043],mul_res1[5044],mul_res1[5045],mul_res1[5046],mul_res1[5047],mul_res1[5048],mul_res1[5049],mul_res1[5050],mul_res1[5051],mul_res1[5052],mul_res1[5053],mul_res1[5054],mul_res1[5055],mul_res1[5056],mul_res1[5057],mul_res1[5058],mul_res1[5059],mul_res1[5060],mul_res1[5061],mul_res1[5062],mul_res1[5063],mul_res1[5064],mul_res1[5065],mul_res1[5066],mul_res1[5067],mul_res1[5068],mul_res1[5069],mul_res1[5070],mul_res1[5071],mul_res1[5072],mul_res1[5073],mul_res1[5074],mul_res1[5075],mul_res1[5076],mul_res1[5077],mul_res1[5078],mul_res1[5079],mul_res1[5080],mul_res1[5081],mul_res1[5082],mul_res1[5083],mul_res1[5084],mul_res1[5085],mul_res1[5086],mul_res1[5087],mul_res1[5088],mul_res1[5089],mul_res1[5090],mul_res1[5091],mul_res1[5092],mul_res1[5093],mul_res1[5094],mul_res1[5095],mul_res1[5096],mul_res1[5097],mul_res1[5098],mul_res1[5099],mul_res1[5100],mul_res1[5101],mul_res1[5102],mul_res1[5103],mul_res1[5104],mul_res1[5105],mul_res1[5106],mul_res1[5107],mul_res1[5108],mul_res1[5109],mul_res1[5110],mul_res1[5111],mul_res1[5112],mul_res1[5113],mul_res1[5114],mul_res1[5115],mul_res1[5116],mul_res1[5117],mul_res1[5118],mul_res1[5119],mul_res1[5120],mul_res1[5121],mul_res1[5122],mul_res1[5123],mul_res1[5124],mul_res1[5125],mul_res1[5126],mul_res1[5127],mul_res1[5128],mul_res1[5129],mul_res1[5130],mul_res1[5131],mul_res1[5132],mul_res1[5133],mul_res1[5134],mul_res1[5135],mul_res1[5136],mul_res1[5137],mul_res1[5138],mul_res1[5139],mul_res1[5140],mul_res1[5141],mul_res1[5142],mul_res1[5143],mul_res1[5144],mul_res1[5145],mul_res1[5146],mul_res1[5147],mul_res1[5148],mul_res1[5149],mul_res1[5150],mul_res1[5151],mul_res1[5152],mul_res1[5153],mul_res1[5154],mul_res1[5155],mul_res1[5156],mul_res1[5157],mul_res1[5158],mul_res1[5159],mul_res1[5160],mul_res1[5161],mul_res1[5162],mul_res1[5163],mul_res1[5164],mul_res1[5165],mul_res1[5166],mul_res1[5167],mul_res1[5168],mul_res1[5169],mul_res1[5170],mul_res1[5171],mul_res1[5172],mul_res1[5173],mul_res1[5174],mul_res1[5175],mul_res1[5176],mul_res1[5177],mul_res1[5178],mul_res1[5179],mul_res1[5180],mul_res1[5181],mul_res1[5182],mul_res1[5183],mul_res1[5184],mul_res1[5185],mul_res1[5186],mul_res1[5187],mul_res1[5188],mul_res1[5189],mul_res1[5190],mul_res1[5191],mul_res1[5192],mul_res1[5193],mul_res1[5194],mul_res1[5195],mul_res1[5196],mul_res1[5197],mul_res1[5198],mul_res1[5199],result_fc1[25]);


adder_200in adder_200in_mod_26(clk,rst,mul_res1[5200],mul_res1[5201],mul_res1[5202],mul_res1[5203],mul_res1[5204],mul_res1[5205],mul_res1[5206],mul_res1[5207],mul_res1[5208],mul_res1[5209],mul_res1[5210],mul_res1[5211],mul_res1[5212],mul_res1[5213],mul_res1[5214],mul_res1[5215],mul_res1[5216],mul_res1[5217],mul_res1[5218],mul_res1[5219],mul_res1[5220],mul_res1[5221],mul_res1[5222],mul_res1[5223],mul_res1[5224],mul_res1[5225],mul_res1[5226],mul_res1[5227],mul_res1[5228],mul_res1[5229],mul_res1[5230],mul_res1[5231],mul_res1[5232],mul_res1[5233],mul_res1[5234],mul_res1[5235],mul_res1[5236],mul_res1[5237],mul_res1[5238],mul_res1[5239],mul_res1[5240],mul_res1[5241],mul_res1[5242],mul_res1[5243],mul_res1[5244],mul_res1[5245],mul_res1[5246],mul_res1[5247],mul_res1[5248],mul_res1[5249],mul_res1[5250],mul_res1[5251],mul_res1[5252],mul_res1[5253],mul_res1[5254],mul_res1[5255],mul_res1[5256],mul_res1[5257],mul_res1[5258],mul_res1[5259],mul_res1[5260],mul_res1[5261],mul_res1[5262],mul_res1[5263],mul_res1[5264],mul_res1[5265],mul_res1[5266],mul_res1[5267],mul_res1[5268],mul_res1[5269],mul_res1[5270],mul_res1[5271],mul_res1[5272],mul_res1[5273],mul_res1[5274],mul_res1[5275],mul_res1[5276],mul_res1[5277],mul_res1[5278],mul_res1[5279],mul_res1[5280],mul_res1[5281],mul_res1[5282],mul_res1[5283],mul_res1[5284],mul_res1[5285],mul_res1[5286],mul_res1[5287],mul_res1[5288],mul_res1[5289],mul_res1[5290],mul_res1[5291],mul_res1[5292],mul_res1[5293],mul_res1[5294],mul_res1[5295],mul_res1[5296],mul_res1[5297],mul_res1[5298],mul_res1[5299],mul_res1[5300],mul_res1[5301],mul_res1[5302],mul_res1[5303],mul_res1[5304],mul_res1[5305],mul_res1[5306],mul_res1[5307],mul_res1[5308],mul_res1[5309],mul_res1[5310],mul_res1[5311],mul_res1[5312],mul_res1[5313],mul_res1[5314],mul_res1[5315],mul_res1[5316],mul_res1[5317],mul_res1[5318],mul_res1[5319],mul_res1[5320],mul_res1[5321],mul_res1[5322],mul_res1[5323],mul_res1[5324],mul_res1[5325],mul_res1[5326],mul_res1[5327],mul_res1[5328],mul_res1[5329],mul_res1[5330],mul_res1[5331],mul_res1[5332],mul_res1[5333],mul_res1[5334],mul_res1[5335],mul_res1[5336],mul_res1[5337],mul_res1[5338],mul_res1[5339],mul_res1[5340],mul_res1[5341],mul_res1[5342],mul_res1[5343],mul_res1[5344],mul_res1[5345],mul_res1[5346],mul_res1[5347],mul_res1[5348],mul_res1[5349],mul_res1[5350],mul_res1[5351],mul_res1[5352],mul_res1[5353],mul_res1[5354],mul_res1[5355],mul_res1[5356],mul_res1[5357],mul_res1[5358],mul_res1[5359],mul_res1[5360],mul_res1[5361],mul_res1[5362],mul_res1[5363],mul_res1[5364],mul_res1[5365],mul_res1[5366],mul_res1[5367],mul_res1[5368],mul_res1[5369],mul_res1[5370],mul_res1[5371],mul_res1[5372],mul_res1[5373],mul_res1[5374],mul_res1[5375],mul_res1[5376],mul_res1[5377],mul_res1[5378],mul_res1[5379],mul_res1[5380],mul_res1[5381],mul_res1[5382],mul_res1[5383],mul_res1[5384],mul_res1[5385],mul_res1[5386],mul_res1[5387],mul_res1[5388],mul_res1[5389],mul_res1[5390],mul_res1[5391],mul_res1[5392],mul_res1[5393],mul_res1[5394],mul_res1[5395],mul_res1[5396],mul_res1[5397],mul_res1[5398],mul_res1[5399],result_fc1[26]);


adder_200in adder_200in_mod_27(clk,rst,mul_res1[5400],mul_res1[5401],mul_res1[5402],mul_res1[5403],mul_res1[5404],mul_res1[5405],mul_res1[5406],mul_res1[5407],mul_res1[5408],mul_res1[5409],mul_res1[5410],mul_res1[5411],mul_res1[5412],mul_res1[5413],mul_res1[5414],mul_res1[5415],mul_res1[5416],mul_res1[5417],mul_res1[5418],mul_res1[5419],mul_res1[5420],mul_res1[5421],mul_res1[5422],mul_res1[5423],mul_res1[5424],mul_res1[5425],mul_res1[5426],mul_res1[5427],mul_res1[5428],mul_res1[5429],mul_res1[5430],mul_res1[5431],mul_res1[5432],mul_res1[5433],mul_res1[5434],mul_res1[5435],mul_res1[5436],mul_res1[5437],mul_res1[5438],mul_res1[5439],mul_res1[5440],mul_res1[5441],mul_res1[5442],mul_res1[5443],mul_res1[5444],mul_res1[5445],mul_res1[5446],mul_res1[5447],mul_res1[5448],mul_res1[5449],mul_res1[5450],mul_res1[5451],mul_res1[5452],mul_res1[5453],mul_res1[5454],mul_res1[5455],mul_res1[5456],mul_res1[5457],mul_res1[5458],mul_res1[5459],mul_res1[5460],mul_res1[5461],mul_res1[5462],mul_res1[5463],mul_res1[5464],mul_res1[5465],mul_res1[5466],mul_res1[5467],mul_res1[5468],mul_res1[5469],mul_res1[5470],mul_res1[5471],mul_res1[5472],mul_res1[5473],mul_res1[5474],mul_res1[5475],mul_res1[5476],mul_res1[5477],mul_res1[5478],mul_res1[5479],mul_res1[5480],mul_res1[5481],mul_res1[5482],mul_res1[5483],mul_res1[5484],mul_res1[5485],mul_res1[5486],mul_res1[5487],mul_res1[5488],mul_res1[5489],mul_res1[5490],mul_res1[5491],mul_res1[5492],mul_res1[5493],mul_res1[5494],mul_res1[5495],mul_res1[5496],mul_res1[5497],mul_res1[5498],mul_res1[5499],mul_res1[5500],mul_res1[5501],mul_res1[5502],mul_res1[5503],mul_res1[5504],mul_res1[5505],mul_res1[5506],mul_res1[5507],mul_res1[5508],mul_res1[5509],mul_res1[5510],mul_res1[5511],mul_res1[5512],mul_res1[5513],mul_res1[5514],mul_res1[5515],mul_res1[5516],mul_res1[5517],mul_res1[5518],mul_res1[5519],mul_res1[5520],mul_res1[5521],mul_res1[5522],mul_res1[5523],mul_res1[5524],mul_res1[5525],mul_res1[5526],mul_res1[5527],mul_res1[5528],mul_res1[5529],mul_res1[5530],mul_res1[5531],mul_res1[5532],mul_res1[5533],mul_res1[5534],mul_res1[5535],mul_res1[5536],mul_res1[5537],mul_res1[5538],mul_res1[5539],mul_res1[5540],mul_res1[5541],mul_res1[5542],mul_res1[5543],mul_res1[5544],mul_res1[5545],mul_res1[5546],mul_res1[5547],mul_res1[5548],mul_res1[5549],mul_res1[5550],mul_res1[5551],mul_res1[5552],mul_res1[5553],mul_res1[5554],mul_res1[5555],mul_res1[5556],mul_res1[5557],mul_res1[5558],mul_res1[5559],mul_res1[5560],mul_res1[5561],mul_res1[5562],mul_res1[5563],mul_res1[5564],mul_res1[5565],mul_res1[5566],mul_res1[5567],mul_res1[5568],mul_res1[5569],mul_res1[5570],mul_res1[5571],mul_res1[5572],mul_res1[5573],mul_res1[5574],mul_res1[5575],mul_res1[5576],mul_res1[5577],mul_res1[5578],mul_res1[5579],mul_res1[5580],mul_res1[5581],mul_res1[5582],mul_res1[5583],mul_res1[5584],mul_res1[5585],mul_res1[5586],mul_res1[5587],mul_res1[5588],mul_res1[5589],mul_res1[5590],mul_res1[5591],mul_res1[5592],mul_res1[5593],mul_res1[5594],mul_res1[5595],mul_res1[5596],mul_res1[5597],mul_res1[5598],mul_res1[5599],result_fc1[27]);


adder_200in adder_200in_mod_28(clk,rst,mul_res1[5600],mul_res1[5601],mul_res1[5602],mul_res1[5603],mul_res1[5604],mul_res1[5605],mul_res1[5606],mul_res1[5607],mul_res1[5608],mul_res1[5609],mul_res1[5610],mul_res1[5611],mul_res1[5612],mul_res1[5613],mul_res1[5614],mul_res1[5615],mul_res1[5616],mul_res1[5617],mul_res1[5618],mul_res1[5619],mul_res1[5620],mul_res1[5621],mul_res1[5622],mul_res1[5623],mul_res1[5624],mul_res1[5625],mul_res1[5626],mul_res1[5627],mul_res1[5628],mul_res1[5629],mul_res1[5630],mul_res1[5631],mul_res1[5632],mul_res1[5633],mul_res1[5634],mul_res1[5635],mul_res1[5636],mul_res1[5637],mul_res1[5638],mul_res1[5639],mul_res1[5640],mul_res1[5641],mul_res1[5642],mul_res1[5643],mul_res1[5644],mul_res1[5645],mul_res1[5646],mul_res1[5647],mul_res1[5648],mul_res1[5649],mul_res1[5650],mul_res1[5651],mul_res1[5652],mul_res1[5653],mul_res1[5654],mul_res1[5655],mul_res1[5656],mul_res1[5657],mul_res1[5658],mul_res1[5659],mul_res1[5660],mul_res1[5661],mul_res1[5662],mul_res1[5663],mul_res1[5664],mul_res1[5665],mul_res1[5666],mul_res1[5667],mul_res1[5668],mul_res1[5669],mul_res1[5670],mul_res1[5671],mul_res1[5672],mul_res1[5673],mul_res1[5674],mul_res1[5675],mul_res1[5676],mul_res1[5677],mul_res1[5678],mul_res1[5679],mul_res1[5680],mul_res1[5681],mul_res1[5682],mul_res1[5683],mul_res1[5684],mul_res1[5685],mul_res1[5686],mul_res1[5687],mul_res1[5688],mul_res1[5689],mul_res1[5690],mul_res1[5691],mul_res1[5692],mul_res1[5693],mul_res1[5694],mul_res1[5695],mul_res1[5696],mul_res1[5697],mul_res1[5698],mul_res1[5699],mul_res1[5700],mul_res1[5701],mul_res1[5702],mul_res1[5703],mul_res1[5704],mul_res1[5705],mul_res1[5706],mul_res1[5707],mul_res1[5708],mul_res1[5709],mul_res1[5710],mul_res1[5711],mul_res1[5712],mul_res1[5713],mul_res1[5714],mul_res1[5715],mul_res1[5716],mul_res1[5717],mul_res1[5718],mul_res1[5719],mul_res1[5720],mul_res1[5721],mul_res1[5722],mul_res1[5723],mul_res1[5724],mul_res1[5725],mul_res1[5726],mul_res1[5727],mul_res1[5728],mul_res1[5729],mul_res1[5730],mul_res1[5731],mul_res1[5732],mul_res1[5733],mul_res1[5734],mul_res1[5735],mul_res1[5736],mul_res1[5737],mul_res1[5738],mul_res1[5739],mul_res1[5740],mul_res1[5741],mul_res1[5742],mul_res1[5743],mul_res1[5744],mul_res1[5745],mul_res1[5746],mul_res1[5747],mul_res1[5748],mul_res1[5749],mul_res1[5750],mul_res1[5751],mul_res1[5752],mul_res1[5753],mul_res1[5754],mul_res1[5755],mul_res1[5756],mul_res1[5757],mul_res1[5758],mul_res1[5759],mul_res1[5760],mul_res1[5761],mul_res1[5762],mul_res1[5763],mul_res1[5764],mul_res1[5765],mul_res1[5766],mul_res1[5767],mul_res1[5768],mul_res1[5769],mul_res1[5770],mul_res1[5771],mul_res1[5772],mul_res1[5773],mul_res1[5774],mul_res1[5775],mul_res1[5776],mul_res1[5777],mul_res1[5778],mul_res1[5779],mul_res1[5780],mul_res1[5781],mul_res1[5782],mul_res1[5783],mul_res1[5784],mul_res1[5785],mul_res1[5786],mul_res1[5787],mul_res1[5788],mul_res1[5789],mul_res1[5790],mul_res1[5791],mul_res1[5792],mul_res1[5793],mul_res1[5794],mul_res1[5795],mul_res1[5796],mul_res1[5797],mul_res1[5798],mul_res1[5799],result_fc1[28]);


adder_200in adder_200in_mod_29(clk,rst,mul_res1[5800],mul_res1[5801],mul_res1[5802],mul_res1[5803],mul_res1[5804],mul_res1[5805],mul_res1[5806],mul_res1[5807],mul_res1[5808],mul_res1[5809],mul_res1[5810],mul_res1[5811],mul_res1[5812],mul_res1[5813],mul_res1[5814],mul_res1[5815],mul_res1[5816],mul_res1[5817],mul_res1[5818],mul_res1[5819],mul_res1[5820],mul_res1[5821],mul_res1[5822],mul_res1[5823],mul_res1[5824],mul_res1[5825],mul_res1[5826],mul_res1[5827],mul_res1[5828],mul_res1[5829],mul_res1[5830],mul_res1[5831],mul_res1[5832],mul_res1[5833],mul_res1[5834],mul_res1[5835],mul_res1[5836],mul_res1[5837],mul_res1[5838],mul_res1[5839],mul_res1[5840],mul_res1[5841],mul_res1[5842],mul_res1[5843],mul_res1[5844],mul_res1[5845],mul_res1[5846],mul_res1[5847],mul_res1[5848],mul_res1[5849],mul_res1[5850],mul_res1[5851],mul_res1[5852],mul_res1[5853],mul_res1[5854],mul_res1[5855],mul_res1[5856],mul_res1[5857],mul_res1[5858],mul_res1[5859],mul_res1[5860],mul_res1[5861],mul_res1[5862],mul_res1[5863],mul_res1[5864],mul_res1[5865],mul_res1[5866],mul_res1[5867],mul_res1[5868],mul_res1[5869],mul_res1[5870],mul_res1[5871],mul_res1[5872],mul_res1[5873],mul_res1[5874],mul_res1[5875],mul_res1[5876],mul_res1[5877],mul_res1[5878],mul_res1[5879],mul_res1[5880],mul_res1[5881],mul_res1[5882],mul_res1[5883],mul_res1[5884],mul_res1[5885],mul_res1[5886],mul_res1[5887],mul_res1[5888],mul_res1[5889],mul_res1[5890],mul_res1[5891],mul_res1[5892],mul_res1[5893],mul_res1[5894],mul_res1[5895],mul_res1[5896],mul_res1[5897],mul_res1[5898],mul_res1[5899],mul_res1[5900],mul_res1[5901],mul_res1[5902],mul_res1[5903],mul_res1[5904],mul_res1[5905],mul_res1[5906],mul_res1[5907],mul_res1[5908],mul_res1[5909],mul_res1[5910],mul_res1[5911],mul_res1[5912],mul_res1[5913],mul_res1[5914],mul_res1[5915],mul_res1[5916],mul_res1[5917],mul_res1[5918],mul_res1[5919],mul_res1[5920],mul_res1[5921],mul_res1[5922],mul_res1[5923],mul_res1[5924],mul_res1[5925],mul_res1[5926],mul_res1[5927],mul_res1[5928],mul_res1[5929],mul_res1[5930],mul_res1[5931],mul_res1[5932],mul_res1[5933],mul_res1[5934],mul_res1[5935],mul_res1[5936],mul_res1[5937],mul_res1[5938],mul_res1[5939],mul_res1[5940],mul_res1[5941],mul_res1[5942],mul_res1[5943],mul_res1[5944],mul_res1[5945],mul_res1[5946],mul_res1[5947],mul_res1[5948],mul_res1[5949],mul_res1[5950],mul_res1[5951],mul_res1[5952],mul_res1[5953],mul_res1[5954],mul_res1[5955],mul_res1[5956],mul_res1[5957],mul_res1[5958],mul_res1[5959],mul_res1[5960],mul_res1[5961],mul_res1[5962],mul_res1[5963],mul_res1[5964],mul_res1[5965],mul_res1[5966],mul_res1[5967],mul_res1[5968],mul_res1[5969],mul_res1[5970],mul_res1[5971],mul_res1[5972],mul_res1[5973],mul_res1[5974],mul_res1[5975],mul_res1[5976],mul_res1[5977],mul_res1[5978],mul_res1[5979],mul_res1[5980],mul_res1[5981],mul_res1[5982],mul_res1[5983],mul_res1[5984],mul_res1[5985],mul_res1[5986],mul_res1[5987],mul_res1[5988],mul_res1[5989],mul_res1[5990],mul_res1[5991],mul_res1[5992],mul_res1[5993],mul_res1[5994],mul_res1[5995],mul_res1[5996],mul_res1[5997],mul_res1[5998],mul_res1[5999],result_fc1[29]);


adder_200in adder_200in_mod_30(clk,rst,mul_res1[6000],mul_res1[6001],mul_res1[6002],mul_res1[6003],mul_res1[6004],mul_res1[6005],mul_res1[6006],mul_res1[6007],mul_res1[6008],mul_res1[6009],mul_res1[6010],mul_res1[6011],mul_res1[6012],mul_res1[6013],mul_res1[6014],mul_res1[6015],mul_res1[6016],mul_res1[6017],mul_res1[6018],mul_res1[6019],mul_res1[6020],mul_res1[6021],mul_res1[6022],mul_res1[6023],mul_res1[6024],mul_res1[6025],mul_res1[6026],mul_res1[6027],mul_res1[6028],mul_res1[6029],mul_res1[6030],mul_res1[6031],mul_res1[6032],mul_res1[6033],mul_res1[6034],mul_res1[6035],mul_res1[6036],mul_res1[6037],mul_res1[6038],mul_res1[6039],mul_res1[6040],mul_res1[6041],mul_res1[6042],mul_res1[6043],mul_res1[6044],mul_res1[6045],mul_res1[6046],mul_res1[6047],mul_res1[6048],mul_res1[6049],mul_res1[6050],mul_res1[6051],mul_res1[6052],mul_res1[6053],mul_res1[6054],mul_res1[6055],mul_res1[6056],mul_res1[6057],mul_res1[6058],mul_res1[6059],mul_res1[6060],mul_res1[6061],mul_res1[6062],mul_res1[6063],mul_res1[6064],mul_res1[6065],mul_res1[6066],mul_res1[6067],mul_res1[6068],mul_res1[6069],mul_res1[6070],mul_res1[6071],mul_res1[6072],mul_res1[6073],mul_res1[6074],mul_res1[6075],mul_res1[6076],mul_res1[6077],mul_res1[6078],mul_res1[6079],mul_res1[6080],mul_res1[6081],mul_res1[6082],mul_res1[6083],mul_res1[6084],mul_res1[6085],mul_res1[6086],mul_res1[6087],mul_res1[6088],mul_res1[6089],mul_res1[6090],mul_res1[6091],mul_res1[6092],mul_res1[6093],mul_res1[6094],mul_res1[6095],mul_res1[6096],mul_res1[6097],mul_res1[6098],mul_res1[6099],mul_res1[6100],mul_res1[6101],mul_res1[6102],mul_res1[6103],mul_res1[6104],mul_res1[6105],mul_res1[6106],mul_res1[6107],mul_res1[6108],mul_res1[6109],mul_res1[6110],mul_res1[6111],mul_res1[6112],mul_res1[6113],mul_res1[6114],mul_res1[6115],mul_res1[6116],mul_res1[6117],mul_res1[6118],mul_res1[6119],mul_res1[6120],mul_res1[6121],mul_res1[6122],mul_res1[6123],mul_res1[6124],mul_res1[6125],mul_res1[6126],mul_res1[6127],mul_res1[6128],mul_res1[6129],mul_res1[6130],mul_res1[6131],mul_res1[6132],mul_res1[6133],mul_res1[6134],mul_res1[6135],mul_res1[6136],mul_res1[6137],mul_res1[6138],mul_res1[6139],mul_res1[6140],mul_res1[6141],mul_res1[6142],mul_res1[6143],mul_res1[6144],mul_res1[6145],mul_res1[6146],mul_res1[6147],mul_res1[6148],mul_res1[6149],mul_res1[6150],mul_res1[6151],mul_res1[6152],mul_res1[6153],mul_res1[6154],mul_res1[6155],mul_res1[6156],mul_res1[6157],mul_res1[6158],mul_res1[6159],mul_res1[6160],mul_res1[6161],mul_res1[6162],mul_res1[6163],mul_res1[6164],mul_res1[6165],mul_res1[6166],mul_res1[6167],mul_res1[6168],mul_res1[6169],mul_res1[6170],mul_res1[6171],mul_res1[6172],mul_res1[6173],mul_res1[6174],mul_res1[6175],mul_res1[6176],mul_res1[6177],mul_res1[6178],mul_res1[6179],mul_res1[6180],mul_res1[6181],mul_res1[6182],mul_res1[6183],mul_res1[6184],mul_res1[6185],mul_res1[6186],mul_res1[6187],mul_res1[6188],mul_res1[6189],mul_res1[6190],mul_res1[6191],mul_res1[6192],mul_res1[6193],mul_res1[6194],mul_res1[6195],mul_res1[6196],mul_res1[6197],mul_res1[6198],mul_res1[6199],result_fc1[30]);


adder_200in adder_200in_mod_31(clk,rst,mul_res1[6200],mul_res1[6201],mul_res1[6202],mul_res1[6203],mul_res1[6204],mul_res1[6205],mul_res1[6206],mul_res1[6207],mul_res1[6208],mul_res1[6209],mul_res1[6210],mul_res1[6211],mul_res1[6212],mul_res1[6213],mul_res1[6214],mul_res1[6215],mul_res1[6216],mul_res1[6217],mul_res1[6218],mul_res1[6219],mul_res1[6220],mul_res1[6221],mul_res1[6222],mul_res1[6223],mul_res1[6224],mul_res1[6225],mul_res1[6226],mul_res1[6227],mul_res1[6228],mul_res1[6229],mul_res1[6230],mul_res1[6231],mul_res1[6232],mul_res1[6233],mul_res1[6234],mul_res1[6235],mul_res1[6236],mul_res1[6237],mul_res1[6238],mul_res1[6239],mul_res1[6240],mul_res1[6241],mul_res1[6242],mul_res1[6243],mul_res1[6244],mul_res1[6245],mul_res1[6246],mul_res1[6247],mul_res1[6248],mul_res1[6249],mul_res1[6250],mul_res1[6251],mul_res1[6252],mul_res1[6253],mul_res1[6254],mul_res1[6255],mul_res1[6256],mul_res1[6257],mul_res1[6258],mul_res1[6259],mul_res1[6260],mul_res1[6261],mul_res1[6262],mul_res1[6263],mul_res1[6264],mul_res1[6265],mul_res1[6266],mul_res1[6267],mul_res1[6268],mul_res1[6269],mul_res1[6270],mul_res1[6271],mul_res1[6272],mul_res1[6273],mul_res1[6274],mul_res1[6275],mul_res1[6276],mul_res1[6277],mul_res1[6278],mul_res1[6279],mul_res1[6280],mul_res1[6281],mul_res1[6282],mul_res1[6283],mul_res1[6284],mul_res1[6285],mul_res1[6286],mul_res1[6287],mul_res1[6288],mul_res1[6289],mul_res1[6290],mul_res1[6291],mul_res1[6292],mul_res1[6293],mul_res1[6294],mul_res1[6295],mul_res1[6296],mul_res1[6297],mul_res1[6298],mul_res1[6299],mul_res1[6300],mul_res1[6301],mul_res1[6302],mul_res1[6303],mul_res1[6304],mul_res1[6305],mul_res1[6306],mul_res1[6307],mul_res1[6308],mul_res1[6309],mul_res1[6310],mul_res1[6311],mul_res1[6312],mul_res1[6313],mul_res1[6314],mul_res1[6315],mul_res1[6316],mul_res1[6317],mul_res1[6318],mul_res1[6319],mul_res1[6320],mul_res1[6321],mul_res1[6322],mul_res1[6323],mul_res1[6324],mul_res1[6325],mul_res1[6326],mul_res1[6327],mul_res1[6328],mul_res1[6329],mul_res1[6330],mul_res1[6331],mul_res1[6332],mul_res1[6333],mul_res1[6334],mul_res1[6335],mul_res1[6336],mul_res1[6337],mul_res1[6338],mul_res1[6339],mul_res1[6340],mul_res1[6341],mul_res1[6342],mul_res1[6343],mul_res1[6344],mul_res1[6345],mul_res1[6346],mul_res1[6347],mul_res1[6348],mul_res1[6349],mul_res1[6350],mul_res1[6351],mul_res1[6352],mul_res1[6353],mul_res1[6354],mul_res1[6355],mul_res1[6356],mul_res1[6357],mul_res1[6358],mul_res1[6359],mul_res1[6360],mul_res1[6361],mul_res1[6362],mul_res1[6363],mul_res1[6364],mul_res1[6365],mul_res1[6366],mul_res1[6367],mul_res1[6368],mul_res1[6369],mul_res1[6370],mul_res1[6371],mul_res1[6372],mul_res1[6373],mul_res1[6374],mul_res1[6375],mul_res1[6376],mul_res1[6377],mul_res1[6378],mul_res1[6379],mul_res1[6380],mul_res1[6381],mul_res1[6382],mul_res1[6383],mul_res1[6384],mul_res1[6385],mul_res1[6386],mul_res1[6387],mul_res1[6388],mul_res1[6389],mul_res1[6390],mul_res1[6391],mul_res1[6392],mul_res1[6393],mul_res1[6394],mul_res1[6395],mul_res1[6396],mul_res1[6397],mul_res1[6398],mul_res1[6399],result_fc1[31]);


adder_200in adder_200in_mod_32(clk,rst,mul_res1[6400],mul_res1[6401],mul_res1[6402],mul_res1[6403],mul_res1[6404],mul_res1[6405],mul_res1[6406],mul_res1[6407],mul_res1[6408],mul_res1[6409],mul_res1[6410],mul_res1[6411],mul_res1[6412],mul_res1[6413],mul_res1[6414],mul_res1[6415],mul_res1[6416],mul_res1[6417],mul_res1[6418],mul_res1[6419],mul_res1[6420],mul_res1[6421],mul_res1[6422],mul_res1[6423],mul_res1[6424],mul_res1[6425],mul_res1[6426],mul_res1[6427],mul_res1[6428],mul_res1[6429],mul_res1[6430],mul_res1[6431],mul_res1[6432],mul_res1[6433],mul_res1[6434],mul_res1[6435],mul_res1[6436],mul_res1[6437],mul_res1[6438],mul_res1[6439],mul_res1[6440],mul_res1[6441],mul_res1[6442],mul_res1[6443],mul_res1[6444],mul_res1[6445],mul_res1[6446],mul_res1[6447],mul_res1[6448],mul_res1[6449],mul_res1[6450],mul_res1[6451],mul_res1[6452],mul_res1[6453],mul_res1[6454],mul_res1[6455],mul_res1[6456],mul_res1[6457],mul_res1[6458],mul_res1[6459],mul_res1[6460],mul_res1[6461],mul_res1[6462],mul_res1[6463],mul_res1[6464],mul_res1[6465],mul_res1[6466],mul_res1[6467],mul_res1[6468],mul_res1[6469],mul_res1[6470],mul_res1[6471],mul_res1[6472],mul_res1[6473],mul_res1[6474],mul_res1[6475],mul_res1[6476],mul_res1[6477],mul_res1[6478],mul_res1[6479],mul_res1[6480],mul_res1[6481],mul_res1[6482],mul_res1[6483],mul_res1[6484],mul_res1[6485],mul_res1[6486],mul_res1[6487],mul_res1[6488],mul_res1[6489],mul_res1[6490],mul_res1[6491],mul_res1[6492],mul_res1[6493],mul_res1[6494],mul_res1[6495],mul_res1[6496],mul_res1[6497],mul_res1[6498],mul_res1[6499],mul_res1[6500],mul_res1[6501],mul_res1[6502],mul_res1[6503],mul_res1[6504],mul_res1[6505],mul_res1[6506],mul_res1[6507],mul_res1[6508],mul_res1[6509],mul_res1[6510],mul_res1[6511],mul_res1[6512],mul_res1[6513],mul_res1[6514],mul_res1[6515],mul_res1[6516],mul_res1[6517],mul_res1[6518],mul_res1[6519],mul_res1[6520],mul_res1[6521],mul_res1[6522],mul_res1[6523],mul_res1[6524],mul_res1[6525],mul_res1[6526],mul_res1[6527],mul_res1[6528],mul_res1[6529],mul_res1[6530],mul_res1[6531],mul_res1[6532],mul_res1[6533],mul_res1[6534],mul_res1[6535],mul_res1[6536],mul_res1[6537],mul_res1[6538],mul_res1[6539],mul_res1[6540],mul_res1[6541],mul_res1[6542],mul_res1[6543],mul_res1[6544],mul_res1[6545],mul_res1[6546],mul_res1[6547],mul_res1[6548],mul_res1[6549],mul_res1[6550],mul_res1[6551],mul_res1[6552],mul_res1[6553],mul_res1[6554],mul_res1[6555],mul_res1[6556],mul_res1[6557],mul_res1[6558],mul_res1[6559],mul_res1[6560],mul_res1[6561],mul_res1[6562],mul_res1[6563],mul_res1[6564],mul_res1[6565],mul_res1[6566],mul_res1[6567],mul_res1[6568],mul_res1[6569],mul_res1[6570],mul_res1[6571],mul_res1[6572],mul_res1[6573],mul_res1[6574],mul_res1[6575],mul_res1[6576],mul_res1[6577],mul_res1[6578],mul_res1[6579],mul_res1[6580],mul_res1[6581],mul_res1[6582],mul_res1[6583],mul_res1[6584],mul_res1[6585],mul_res1[6586],mul_res1[6587],mul_res1[6588],mul_res1[6589],mul_res1[6590],mul_res1[6591],mul_res1[6592],mul_res1[6593],mul_res1[6594],mul_res1[6595],mul_res1[6596],mul_res1[6597],mul_res1[6598],mul_res1[6599],result_fc1[32]);


adder_200in adder_200in_mod_33(clk,rst,mul_res1[6600],mul_res1[6601],mul_res1[6602],mul_res1[6603],mul_res1[6604],mul_res1[6605],mul_res1[6606],mul_res1[6607],mul_res1[6608],mul_res1[6609],mul_res1[6610],mul_res1[6611],mul_res1[6612],mul_res1[6613],mul_res1[6614],mul_res1[6615],mul_res1[6616],mul_res1[6617],mul_res1[6618],mul_res1[6619],mul_res1[6620],mul_res1[6621],mul_res1[6622],mul_res1[6623],mul_res1[6624],mul_res1[6625],mul_res1[6626],mul_res1[6627],mul_res1[6628],mul_res1[6629],mul_res1[6630],mul_res1[6631],mul_res1[6632],mul_res1[6633],mul_res1[6634],mul_res1[6635],mul_res1[6636],mul_res1[6637],mul_res1[6638],mul_res1[6639],mul_res1[6640],mul_res1[6641],mul_res1[6642],mul_res1[6643],mul_res1[6644],mul_res1[6645],mul_res1[6646],mul_res1[6647],mul_res1[6648],mul_res1[6649],mul_res1[6650],mul_res1[6651],mul_res1[6652],mul_res1[6653],mul_res1[6654],mul_res1[6655],mul_res1[6656],mul_res1[6657],mul_res1[6658],mul_res1[6659],mul_res1[6660],mul_res1[6661],mul_res1[6662],mul_res1[6663],mul_res1[6664],mul_res1[6665],mul_res1[6666],mul_res1[6667],mul_res1[6668],mul_res1[6669],mul_res1[6670],mul_res1[6671],mul_res1[6672],mul_res1[6673],mul_res1[6674],mul_res1[6675],mul_res1[6676],mul_res1[6677],mul_res1[6678],mul_res1[6679],mul_res1[6680],mul_res1[6681],mul_res1[6682],mul_res1[6683],mul_res1[6684],mul_res1[6685],mul_res1[6686],mul_res1[6687],mul_res1[6688],mul_res1[6689],mul_res1[6690],mul_res1[6691],mul_res1[6692],mul_res1[6693],mul_res1[6694],mul_res1[6695],mul_res1[6696],mul_res1[6697],mul_res1[6698],mul_res1[6699],mul_res1[6700],mul_res1[6701],mul_res1[6702],mul_res1[6703],mul_res1[6704],mul_res1[6705],mul_res1[6706],mul_res1[6707],mul_res1[6708],mul_res1[6709],mul_res1[6710],mul_res1[6711],mul_res1[6712],mul_res1[6713],mul_res1[6714],mul_res1[6715],mul_res1[6716],mul_res1[6717],mul_res1[6718],mul_res1[6719],mul_res1[6720],mul_res1[6721],mul_res1[6722],mul_res1[6723],mul_res1[6724],mul_res1[6725],mul_res1[6726],mul_res1[6727],mul_res1[6728],mul_res1[6729],mul_res1[6730],mul_res1[6731],mul_res1[6732],mul_res1[6733],mul_res1[6734],mul_res1[6735],mul_res1[6736],mul_res1[6737],mul_res1[6738],mul_res1[6739],mul_res1[6740],mul_res1[6741],mul_res1[6742],mul_res1[6743],mul_res1[6744],mul_res1[6745],mul_res1[6746],mul_res1[6747],mul_res1[6748],mul_res1[6749],mul_res1[6750],mul_res1[6751],mul_res1[6752],mul_res1[6753],mul_res1[6754],mul_res1[6755],mul_res1[6756],mul_res1[6757],mul_res1[6758],mul_res1[6759],mul_res1[6760],mul_res1[6761],mul_res1[6762],mul_res1[6763],mul_res1[6764],mul_res1[6765],mul_res1[6766],mul_res1[6767],mul_res1[6768],mul_res1[6769],mul_res1[6770],mul_res1[6771],mul_res1[6772],mul_res1[6773],mul_res1[6774],mul_res1[6775],mul_res1[6776],mul_res1[6777],mul_res1[6778],mul_res1[6779],mul_res1[6780],mul_res1[6781],mul_res1[6782],mul_res1[6783],mul_res1[6784],mul_res1[6785],mul_res1[6786],mul_res1[6787],mul_res1[6788],mul_res1[6789],mul_res1[6790],mul_res1[6791],mul_res1[6792],mul_res1[6793],mul_res1[6794],mul_res1[6795],mul_res1[6796],mul_res1[6797],mul_res1[6798],mul_res1[6799],result_fc1[33]);


adder_200in adder_200in_mod_34(clk,rst,mul_res1[6800],mul_res1[6801],mul_res1[6802],mul_res1[6803],mul_res1[6804],mul_res1[6805],mul_res1[6806],mul_res1[6807],mul_res1[6808],mul_res1[6809],mul_res1[6810],mul_res1[6811],mul_res1[6812],mul_res1[6813],mul_res1[6814],mul_res1[6815],mul_res1[6816],mul_res1[6817],mul_res1[6818],mul_res1[6819],mul_res1[6820],mul_res1[6821],mul_res1[6822],mul_res1[6823],mul_res1[6824],mul_res1[6825],mul_res1[6826],mul_res1[6827],mul_res1[6828],mul_res1[6829],mul_res1[6830],mul_res1[6831],mul_res1[6832],mul_res1[6833],mul_res1[6834],mul_res1[6835],mul_res1[6836],mul_res1[6837],mul_res1[6838],mul_res1[6839],mul_res1[6840],mul_res1[6841],mul_res1[6842],mul_res1[6843],mul_res1[6844],mul_res1[6845],mul_res1[6846],mul_res1[6847],mul_res1[6848],mul_res1[6849],mul_res1[6850],mul_res1[6851],mul_res1[6852],mul_res1[6853],mul_res1[6854],mul_res1[6855],mul_res1[6856],mul_res1[6857],mul_res1[6858],mul_res1[6859],mul_res1[6860],mul_res1[6861],mul_res1[6862],mul_res1[6863],mul_res1[6864],mul_res1[6865],mul_res1[6866],mul_res1[6867],mul_res1[6868],mul_res1[6869],mul_res1[6870],mul_res1[6871],mul_res1[6872],mul_res1[6873],mul_res1[6874],mul_res1[6875],mul_res1[6876],mul_res1[6877],mul_res1[6878],mul_res1[6879],mul_res1[6880],mul_res1[6881],mul_res1[6882],mul_res1[6883],mul_res1[6884],mul_res1[6885],mul_res1[6886],mul_res1[6887],mul_res1[6888],mul_res1[6889],mul_res1[6890],mul_res1[6891],mul_res1[6892],mul_res1[6893],mul_res1[6894],mul_res1[6895],mul_res1[6896],mul_res1[6897],mul_res1[6898],mul_res1[6899],mul_res1[6900],mul_res1[6901],mul_res1[6902],mul_res1[6903],mul_res1[6904],mul_res1[6905],mul_res1[6906],mul_res1[6907],mul_res1[6908],mul_res1[6909],mul_res1[6910],mul_res1[6911],mul_res1[6912],mul_res1[6913],mul_res1[6914],mul_res1[6915],mul_res1[6916],mul_res1[6917],mul_res1[6918],mul_res1[6919],mul_res1[6920],mul_res1[6921],mul_res1[6922],mul_res1[6923],mul_res1[6924],mul_res1[6925],mul_res1[6926],mul_res1[6927],mul_res1[6928],mul_res1[6929],mul_res1[6930],mul_res1[6931],mul_res1[6932],mul_res1[6933],mul_res1[6934],mul_res1[6935],mul_res1[6936],mul_res1[6937],mul_res1[6938],mul_res1[6939],mul_res1[6940],mul_res1[6941],mul_res1[6942],mul_res1[6943],mul_res1[6944],mul_res1[6945],mul_res1[6946],mul_res1[6947],mul_res1[6948],mul_res1[6949],mul_res1[6950],mul_res1[6951],mul_res1[6952],mul_res1[6953],mul_res1[6954],mul_res1[6955],mul_res1[6956],mul_res1[6957],mul_res1[6958],mul_res1[6959],mul_res1[6960],mul_res1[6961],mul_res1[6962],mul_res1[6963],mul_res1[6964],mul_res1[6965],mul_res1[6966],mul_res1[6967],mul_res1[6968],mul_res1[6969],mul_res1[6970],mul_res1[6971],mul_res1[6972],mul_res1[6973],mul_res1[6974],mul_res1[6975],mul_res1[6976],mul_res1[6977],mul_res1[6978],mul_res1[6979],mul_res1[6980],mul_res1[6981],mul_res1[6982],mul_res1[6983],mul_res1[6984],mul_res1[6985],mul_res1[6986],mul_res1[6987],mul_res1[6988],mul_res1[6989],mul_res1[6990],mul_res1[6991],mul_res1[6992],mul_res1[6993],mul_res1[6994],mul_res1[6995],mul_res1[6996],mul_res1[6997],mul_res1[6998],mul_res1[6999],result_fc1[34]);


adder_200in adder_200in_mod_35(clk,rst,mul_res1[7000],mul_res1[7001],mul_res1[7002],mul_res1[7003],mul_res1[7004],mul_res1[7005],mul_res1[7006],mul_res1[7007],mul_res1[7008],mul_res1[7009],mul_res1[7010],mul_res1[7011],mul_res1[7012],mul_res1[7013],mul_res1[7014],mul_res1[7015],mul_res1[7016],mul_res1[7017],mul_res1[7018],mul_res1[7019],mul_res1[7020],mul_res1[7021],mul_res1[7022],mul_res1[7023],mul_res1[7024],mul_res1[7025],mul_res1[7026],mul_res1[7027],mul_res1[7028],mul_res1[7029],mul_res1[7030],mul_res1[7031],mul_res1[7032],mul_res1[7033],mul_res1[7034],mul_res1[7035],mul_res1[7036],mul_res1[7037],mul_res1[7038],mul_res1[7039],mul_res1[7040],mul_res1[7041],mul_res1[7042],mul_res1[7043],mul_res1[7044],mul_res1[7045],mul_res1[7046],mul_res1[7047],mul_res1[7048],mul_res1[7049],mul_res1[7050],mul_res1[7051],mul_res1[7052],mul_res1[7053],mul_res1[7054],mul_res1[7055],mul_res1[7056],mul_res1[7057],mul_res1[7058],mul_res1[7059],mul_res1[7060],mul_res1[7061],mul_res1[7062],mul_res1[7063],mul_res1[7064],mul_res1[7065],mul_res1[7066],mul_res1[7067],mul_res1[7068],mul_res1[7069],mul_res1[7070],mul_res1[7071],mul_res1[7072],mul_res1[7073],mul_res1[7074],mul_res1[7075],mul_res1[7076],mul_res1[7077],mul_res1[7078],mul_res1[7079],mul_res1[7080],mul_res1[7081],mul_res1[7082],mul_res1[7083],mul_res1[7084],mul_res1[7085],mul_res1[7086],mul_res1[7087],mul_res1[7088],mul_res1[7089],mul_res1[7090],mul_res1[7091],mul_res1[7092],mul_res1[7093],mul_res1[7094],mul_res1[7095],mul_res1[7096],mul_res1[7097],mul_res1[7098],mul_res1[7099],mul_res1[7100],mul_res1[7101],mul_res1[7102],mul_res1[7103],mul_res1[7104],mul_res1[7105],mul_res1[7106],mul_res1[7107],mul_res1[7108],mul_res1[7109],mul_res1[7110],mul_res1[7111],mul_res1[7112],mul_res1[7113],mul_res1[7114],mul_res1[7115],mul_res1[7116],mul_res1[7117],mul_res1[7118],mul_res1[7119],mul_res1[7120],mul_res1[7121],mul_res1[7122],mul_res1[7123],mul_res1[7124],mul_res1[7125],mul_res1[7126],mul_res1[7127],mul_res1[7128],mul_res1[7129],mul_res1[7130],mul_res1[7131],mul_res1[7132],mul_res1[7133],mul_res1[7134],mul_res1[7135],mul_res1[7136],mul_res1[7137],mul_res1[7138],mul_res1[7139],mul_res1[7140],mul_res1[7141],mul_res1[7142],mul_res1[7143],mul_res1[7144],mul_res1[7145],mul_res1[7146],mul_res1[7147],mul_res1[7148],mul_res1[7149],mul_res1[7150],mul_res1[7151],mul_res1[7152],mul_res1[7153],mul_res1[7154],mul_res1[7155],mul_res1[7156],mul_res1[7157],mul_res1[7158],mul_res1[7159],mul_res1[7160],mul_res1[7161],mul_res1[7162],mul_res1[7163],mul_res1[7164],mul_res1[7165],mul_res1[7166],mul_res1[7167],mul_res1[7168],mul_res1[7169],mul_res1[7170],mul_res1[7171],mul_res1[7172],mul_res1[7173],mul_res1[7174],mul_res1[7175],mul_res1[7176],mul_res1[7177],mul_res1[7178],mul_res1[7179],mul_res1[7180],mul_res1[7181],mul_res1[7182],mul_res1[7183],mul_res1[7184],mul_res1[7185],mul_res1[7186],mul_res1[7187],mul_res1[7188],mul_res1[7189],mul_res1[7190],mul_res1[7191],mul_res1[7192],mul_res1[7193],mul_res1[7194],mul_res1[7195],mul_res1[7196],mul_res1[7197],mul_res1[7198],mul_res1[7199],result_fc1[35]);


adder_200in adder_200in_mod_36(clk,rst,mul_res1[7200],mul_res1[7201],mul_res1[7202],mul_res1[7203],mul_res1[7204],mul_res1[7205],mul_res1[7206],mul_res1[7207],mul_res1[7208],mul_res1[7209],mul_res1[7210],mul_res1[7211],mul_res1[7212],mul_res1[7213],mul_res1[7214],mul_res1[7215],mul_res1[7216],mul_res1[7217],mul_res1[7218],mul_res1[7219],mul_res1[7220],mul_res1[7221],mul_res1[7222],mul_res1[7223],mul_res1[7224],mul_res1[7225],mul_res1[7226],mul_res1[7227],mul_res1[7228],mul_res1[7229],mul_res1[7230],mul_res1[7231],mul_res1[7232],mul_res1[7233],mul_res1[7234],mul_res1[7235],mul_res1[7236],mul_res1[7237],mul_res1[7238],mul_res1[7239],mul_res1[7240],mul_res1[7241],mul_res1[7242],mul_res1[7243],mul_res1[7244],mul_res1[7245],mul_res1[7246],mul_res1[7247],mul_res1[7248],mul_res1[7249],mul_res1[7250],mul_res1[7251],mul_res1[7252],mul_res1[7253],mul_res1[7254],mul_res1[7255],mul_res1[7256],mul_res1[7257],mul_res1[7258],mul_res1[7259],mul_res1[7260],mul_res1[7261],mul_res1[7262],mul_res1[7263],mul_res1[7264],mul_res1[7265],mul_res1[7266],mul_res1[7267],mul_res1[7268],mul_res1[7269],mul_res1[7270],mul_res1[7271],mul_res1[7272],mul_res1[7273],mul_res1[7274],mul_res1[7275],mul_res1[7276],mul_res1[7277],mul_res1[7278],mul_res1[7279],mul_res1[7280],mul_res1[7281],mul_res1[7282],mul_res1[7283],mul_res1[7284],mul_res1[7285],mul_res1[7286],mul_res1[7287],mul_res1[7288],mul_res1[7289],mul_res1[7290],mul_res1[7291],mul_res1[7292],mul_res1[7293],mul_res1[7294],mul_res1[7295],mul_res1[7296],mul_res1[7297],mul_res1[7298],mul_res1[7299],mul_res1[7300],mul_res1[7301],mul_res1[7302],mul_res1[7303],mul_res1[7304],mul_res1[7305],mul_res1[7306],mul_res1[7307],mul_res1[7308],mul_res1[7309],mul_res1[7310],mul_res1[7311],mul_res1[7312],mul_res1[7313],mul_res1[7314],mul_res1[7315],mul_res1[7316],mul_res1[7317],mul_res1[7318],mul_res1[7319],mul_res1[7320],mul_res1[7321],mul_res1[7322],mul_res1[7323],mul_res1[7324],mul_res1[7325],mul_res1[7326],mul_res1[7327],mul_res1[7328],mul_res1[7329],mul_res1[7330],mul_res1[7331],mul_res1[7332],mul_res1[7333],mul_res1[7334],mul_res1[7335],mul_res1[7336],mul_res1[7337],mul_res1[7338],mul_res1[7339],mul_res1[7340],mul_res1[7341],mul_res1[7342],mul_res1[7343],mul_res1[7344],mul_res1[7345],mul_res1[7346],mul_res1[7347],mul_res1[7348],mul_res1[7349],mul_res1[7350],mul_res1[7351],mul_res1[7352],mul_res1[7353],mul_res1[7354],mul_res1[7355],mul_res1[7356],mul_res1[7357],mul_res1[7358],mul_res1[7359],mul_res1[7360],mul_res1[7361],mul_res1[7362],mul_res1[7363],mul_res1[7364],mul_res1[7365],mul_res1[7366],mul_res1[7367],mul_res1[7368],mul_res1[7369],mul_res1[7370],mul_res1[7371],mul_res1[7372],mul_res1[7373],mul_res1[7374],mul_res1[7375],mul_res1[7376],mul_res1[7377],mul_res1[7378],mul_res1[7379],mul_res1[7380],mul_res1[7381],mul_res1[7382],mul_res1[7383],mul_res1[7384],mul_res1[7385],mul_res1[7386],mul_res1[7387],mul_res1[7388],mul_res1[7389],mul_res1[7390],mul_res1[7391],mul_res1[7392],mul_res1[7393],mul_res1[7394],mul_res1[7395],mul_res1[7396],mul_res1[7397],mul_res1[7398],mul_res1[7399],result_fc1[36]);


adder_200in adder_200in_mod_37(clk,rst,mul_res1[7400],mul_res1[7401],mul_res1[7402],mul_res1[7403],mul_res1[7404],mul_res1[7405],mul_res1[7406],mul_res1[7407],mul_res1[7408],mul_res1[7409],mul_res1[7410],mul_res1[7411],mul_res1[7412],mul_res1[7413],mul_res1[7414],mul_res1[7415],mul_res1[7416],mul_res1[7417],mul_res1[7418],mul_res1[7419],mul_res1[7420],mul_res1[7421],mul_res1[7422],mul_res1[7423],mul_res1[7424],mul_res1[7425],mul_res1[7426],mul_res1[7427],mul_res1[7428],mul_res1[7429],mul_res1[7430],mul_res1[7431],mul_res1[7432],mul_res1[7433],mul_res1[7434],mul_res1[7435],mul_res1[7436],mul_res1[7437],mul_res1[7438],mul_res1[7439],mul_res1[7440],mul_res1[7441],mul_res1[7442],mul_res1[7443],mul_res1[7444],mul_res1[7445],mul_res1[7446],mul_res1[7447],mul_res1[7448],mul_res1[7449],mul_res1[7450],mul_res1[7451],mul_res1[7452],mul_res1[7453],mul_res1[7454],mul_res1[7455],mul_res1[7456],mul_res1[7457],mul_res1[7458],mul_res1[7459],mul_res1[7460],mul_res1[7461],mul_res1[7462],mul_res1[7463],mul_res1[7464],mul_res1[7465],mul_res1[7466],mul_res1[7467],mul_res1[7468],mul_res1[7469],mul_res1[7470],mul_res1[7471],mul_res1[7472],mul_res1[7473],mul_res1[7474],mul_res1[7475],mul_res1[7476],mul_res1[7477],mul_res1[7478],mul_res1[7479],mul_res1[7480],mul_res1[7481],mul_res1[7482],mul_res1[7483],mul_res1[7484],mul_res1[7485],mul_res1[7486],mul_res1[7487],mul_res1[7488],mul_res1[7489],mul_res1[7490],mul_res1[7491],mul_res1[7492],mul_res1[7493],mul_res1[7494],mul_res1[7495],mul_res1[7496],mul_res1[7497],mul_res1[7498],mul_res1[7499],mul_res1[7500],mul_res1[7501],mul_res1[7502],mul_res1[7503],mul_res1[7504],mul_res1[7505],mul_res1[7506],mul_res1[7507],mul_res1[7508],mul_res1[7509],mul_res1[7510],mul_res1[7511],mul_res1[7512],mul_res1[7513],mul_res1[7514],mul_res1[7515],mul_res1[7516],mul_res1[7517],mul_res1[7518],mul_res1[7519],mul_res1[7520],mul_res1[7521],mul_res1[7522],mul_res1[7523],mul_res1[7524],mul_res1[7525],mul_res1[7526],mul_res1[7527],mul_res1[7528],mul_res1[7529],mul_res1[7530],mul_res1[7531],mul_res1[7532],mul_res1[7533],mul_res1[7534],mul_res1[7535],mul_res1[7536],mul_res1[7537],mul_res1[7538],mul_res1[7539],mul_res1[7540],mul_res1[7541],mul_res1[7542],mul_res1[7543],mul_res1[7544],mul_res1[7545],mul_res1[7546],mul_res1[7547],mul_res1[7548],mul_res1[7549],mul_res1[7550],mul_res1[7551],mul_res1[7552],mul_res1[7553],mul_res1[7554],mul_res1[7555],mul_res1[7556],mul_res1[7557],mul_res1[7558],mul_res1[7559],mul_res1[7560],mul_res1[7561],mul_res1[7562],mul_res1[7563],mul_res1[7564],mul_res1[7565],mul_res1[7566],mul_res1[7567],mul_res1[7568],mul_res1[7569],mul_res1[7570],mul_res1[7571],mul_res1[7572],mul_res1[7573],mul_res1[7574],mul_res1[7575],mul_res1[7576],mul_res1[7577],mul_res1[7578],mul_res1[7579],mul_res1[7580],mul_res1[7581],mul_res1[7582],mul_res1[7583],mul_res1[7584],mul_res1[7585],mul_res1[7586],mul_res1[7587],mul_res1[7588],mul_res1[7589],mul_res1[7590],mul_res1[7591],mul_res1[7592],mul_res1[7593],mul_res1[7594],mul_res1[7595],mul_res1[7596],mul_res1[7597],mul_res1[7598],mul_res1[7599],result_fc1[37]);


adder_200in adder_200in_mod_38(clk,rst,mul_res1[7600],mul_res1[7601],mul_res1[7602],mul_res1[7603],mul_res1[7604],mul_res1[7605],mul_res1[7606],mul_res1[7607],mul_res1[7608],mul_res1[7609],mul_res1[7610],mul_res1[7611],mul_res1[7612],mul_res1[7613],mul_res1[7614],mul_res1[7615],mul_res1[7616],mul_res1[7617],mul_res1[7618],mul_res1[7619],mul_res1[7620],mul_res1[7621],mul_res1[7622],mul_res1[7623],mul_res1[7624],mul_res1[7625],mul_res1[7626],mul_res1[7627],mul_res1[7628],mul_res1[7629],mul_res1[7630],mul_res1[7631],mul_res1[7632],mul_res1[7633],mul_res1[7634],mul_res1[7635],mul_res1[7636],mul_res1[7637],mul_res1[7638],mul_res1[7639],mul_res1[7640],mul_res1[7641],mul_res1[7642],mul_res1[7643],mul_res1[7644],mul_res1[7645],mul_res1[7646],mul_res1[7647],mul_res1[7648],mul_res1[7649],mul_res1[7650],mul_res1[7651],mul_res1[7652],mul_res1[7653],mul_res1[7654],mul_res1[7655],mul_res1[7656],mul_res1[7657],mul_res1[7658],mul_res1[7659],mul_res1[7660],mul_res1[7661],mul_res1[7662],mul_res1[7663],mul_res1[7664],mul_res1[7665],mul_res1[7666],mul_res1[7667],mul_res1[7668],mul_res1[7669],mul_res1[7670],mul_res1[7671],mul_res1[7672],mul_res1[7673],mul_res1[7674],mul_res1[7675],mul_res1[7676],mul_res1[7677],mul_res1[7678],mul_res1[7679],mul_res1[7680],mul_res1[7681],mul_res1[7682],mul_res1[7683],mul_res1[7684],mul_res1[7685],mul_res1[7686],mul_res1[7687],mul_res1[7688],mul_res1[7689],mul_res1[7690],mul_res1[7691],mul_res1[7692],mul_res1[7693],mul_res1[7694],mul_res1[7695],mul_res1[7696],mul_res1[7697],mul_res1[7698],mul_res1[7699],mul_res1[7700],mul_res1[7701],mul_res1[7702],mul_res1[7703],mul_res1[7704],mul_res1[7705],mul_res1[7706],mul_res1[7707],mul_res1[7708],mul_res1[7709],mul_res1[7710],mul_res1[7711],mul_res1[7712],mul_res1[7713],mul_res1[7714],mul_res1[7715],mul_res1[7716],mul_res1[7717],mul_res1[7718],mul_res1[7719],mul_res1[7720],mul_res1[7721],mul_res1[7722],mul_res1[7723],mul_res1[7724],mul_res1[7725],mul_res1[7726],mul_res1[7727],mul_res1[7728],mul_res1[7729],mul_res1[7730],mul_res1[7731],mul_res1[7732],mul_res1[7733],mul_res1[7734],mul_res1[7735],mul_res1[7736],mul_res1[7737],mul_res1[7738],mul_res1[7739],mul_res1[7740],mul_res1[7741],mul_res1[7742],mul_res1[7743],mul_res1[7744],mul_res1[7745],mul_res1[7746],mul_res1[7747],mul_res1[7748],mul_res1[7749],mul_res1[7750],mul_res1[7751],mul_res1[7752],mul_res1[7753],mul_res1[7754],mul_res1[7755],mul_res1[7756],mul_res1[7757],mul_res1[7758],mul_res1[7759],mul_res1[7760],mul_res1[7761],mul_res1[7762],mul_res1[7763],mul_res1[7764],mul_res1[7765],mul_res1[7766],mul_res1[7767],mul_res1[7768],mul_res1[7769],mul_res1[7770],mul_res1[7771],mul_res1[7772],mul_res1[7773],mul_res1[7774],mul_res1[7775],mul_res1[7776],mul_res1[7777],mul_res1[7778],mul_res1[7779],mul_res1[7780],mul_res1[7781],mul_res1[7782],mul_res1[7783],mul_res1[7784],mul_res1[7785],mul_res1[7786],mul_res1[7787],mul_res1[7788],mul_res1[7789],mul_res1[7790],mul_res1[7791],mul_res1[7792],mul_res1[7793],mul_res1[7794],mul_res1[7795],mul_res1[7796],mul_res1[7797],mul_res1[7798],mul_res1[7799],result_fc1[38]);


adder_200in adder_200in_mod_39(clk,rst,mul_res1[7800],mul_res1[7801],mul_res1[7802],mul_res1[7803],mul_res1[7804],mul_res1[7805],mul_res1[7806],mul_res1[7807],mul_res1[7808],mul_res1[7809],mul_res1[7810],mul_res1[7811],mul_res1[7812],mul_res1[7813],mul_res1[7814],mul_res1[7815],mul_res1[7816],mul_res1[7817],mul_res1[7818],mul_res1[7819],mul_res1[7820],mul_res1[7821],mul_res1[7822],mul_res1[7823],mul_res1[7824],mul_res1[7825],mul_res1[7826],mul_res1[7827],mul_res1[7828],mul_res1[7829],mul_res1[7830],mul_res1[7831],mul_res1[7832],mul_res1[7833],mul_res1[7834],mul_res1[7835],mul_res1[7836],mul_res1[7837],mul_res1[7838],mul_res1[7839],mul_res1[7840],mul_res1[7841],mul_res1[7842],mul_res1[7843],mul_res1[7844],mul_res1[7845],mul_res1[7846],mul_res1[7847],mul_res1[7848],mul_res1[7849],mul_res1[7850],mul_res1[7851],mul_res1[7852],mul_res1[7853],mul_res1[7854],mul_res1[7855],mul_res1[7856],mul_res1[7857],mul_res1[7858],mul_res1[7859],mul_res1[7860],mul_res1[7861],mul_res1[7862],mul_res1[7863],mul_res1[7864],mul_res1[7865],mul_res1[7866],mul_res1[7867],mul_res1[7868],mul_res1[7869],mul_res1[7870],mul_res1[7871],mul_res1[7872],mul_res1[7873],mul_res1[7874],mul_res1[7875],mul_res1[7876],mul_res1[7877],mul_res1[7878],mul_res1[7879],mul_res1[7880],mul_res1[7881],mul_res1[7882],mul_res1[7883],mul_res1[7884],mul_res1[7885],mul_res1[7886],mul_res1[7887],mul_res1[7888],mul_res1[7889],mul_res1[7890],mul_res1[7891],mul_res1[7892],mul_res1[7893],mul_res1[7894],mul_res1[7895],mul_res1[7896],mul_res1[7897],mul_res1[7898],mul_res1[7899],mul_res1[7900],mul_res1[7901],mul_res1[7902],mul_res1[7903],mul_res1[7904],mul_res1[7905],mul_res1[7906],mul_res1[7907],mul_res1[7908],mul_res1[7909],mul_res1[7910],mul_res1[7911],mul_res1[7912],mul_res1[7913],mul_res1[7914],mul_res1[7915],mul_res1[7916],mul_res1[7917],mul_res1[7918],mul_res1[7919],mul_res1[7920],mul_res1[7921],mul_res1[7922],mul_res1[7923],mul_res1[7924],mul_res1[7925],mul_res1[7926],mul_res1[7927],mul_res1[7928],mul_res1[7929],mul_res1[7930],mul_res1[7931],mul_res1[7932],mul_res1[7933],mul_res1[7934],mul_res1[7935],mul_res1[7936],mul_res1[7937],mul_res1[7938],mul_res1[7939],mul_res1[7940],mul_res1[7941],mul_res1[7942],mul_res1[7943],mul_res1[7944],mul_res1[7945],mul_res1[7946],mul_res1[7947],mul_res1[7948],mul_res1[7949],mul_res1[7950],mul_res1[7951],mul_res1[7952],mul_res1[7953],mul_res1[7954],mul_res1[7955],mul_res1[7956],mul_res1[7957],mul_res1[7958],mul_res1[7959],mul_res1[7960],mul_res1[7961],mul_res1[7962],mul_res1[7963],mul_res1[7964],mul_res1[7965],mul_res1[7966],mul_res1[7967],mul_res1[7968],mul_res1[7969],mul_res1[7970],mul_res1[7971],mul_res1[7972],mul_res1[7973],mul_res1[7974],mul_res1[7975],mul_res1[7976],mul_res1[7977],mul_res1[7978],mul_res1[7979],mul_res1[7980],mul_res1[7981],mul_res1[7982],mul_res1[7983],mul_res1[7984],mul_res1[7985],mul_res1[7986],mul_res1[7987],mul_res1[7988],mul_res1[7989],mul_res1[7990],mul_res1[7991],mul_res1[7992],mul_res1[7993],mul_res1[7994],mul_res1[7995],mul_res1[7996],mul_res1[7997],mul_res1[7998],mul_res1[7999],result_fc1[39]);


adder_200in adder_200in_mod_40(clk,rst,mul_res1[8000],mul_res1[8001],mul_res1[8002],mul_res1[8003],mul_res1[8004],mul_res1[8005],mul_res1[8006],mul_res1[8007],mul_res1[8008],mul_res1[8009],mul_res1[8010],mul_res1[8011],mul_res1[8012],mul_res1[8013],mul_res1[8014],mul_res1[8015],mul_res1[8016],mul_res1[8017],mul_res1[8018],mul_res1[8019],mul_res1[8020],mul_res1[8021],mul_res1[8022],mul_res1[8023],mul_res1[8024],mul_res1[8025],mul_res1[8026],mul_res1[8027],mul_res1[8028],mul_res1[8029],mul_res1[8030],mul_res1[8031],mul_res1[8032],mul_res1[8033],mul_res1[8034],mul_res1[8035],mul_res1[8036],mul_res1[8037],mul_res1[8038],mul_res1[8039],mul_res1[8040],mul_res1[8041],mul_res1[8042],mul_res1[8043],mul_res1[8044],mul_res1[8045],mul_res1[8046],mul_res1[8047],mul_res1[8048],mul_res1[8049],mul_res1[8050],mul_res1[8051],mul_res1[8052],mul_res1[8053],mul_res1[8054],mul_res1[8055],mul_res1[8056],mul_res1[8057],mul_res1[8058],mul_res1[8059],mul_res1[8060],mul_res1[8061],mul_res1[8062],mul_res1[8063],mul_res1[8064],mul_res1[8065],mul_res1[8066],mul_res1[8067],mul_res1[8068],mul_res1[8069],mul_res1[8070],mul_res1[8071],mul_res1[8072],mul_res1[8073],mul_res1[8074],mul_res1[8075],mul_res1[8076],mul_res1[8077],mul_res1[8078],mul_res1[8079],mul_res1[8080],mul_res1[8081],mul_res1[8082],mul_res1[8083],mul_res1[8084],mul_res1[8085],mul_res1[8086],mul_res1[8087],mul_res1[8088],mul_res1[8089],mul_res1[8090],mul_res1[8091],mul_res1[8092],mul_res1[8093],mul_res1[8094],mul_res1[8095],mul_res1[8096],mul_res1[8097],mul_res1[8098],mul_res1[8099],mul_res1[8100],mul_res1[8101],mul_res1[8102],mul_res1[8103],mul_res1[8104],mul_res1[8105],mul_res1[8106],mul_res1[8107],mul_res1[8108],mul_res1[8109],mul_res1[8110],mul_res1[8111],mul_res1[8112],mul_res1[8113],mul_res1[8114],mul_res1[8115],mul_res1[8116],mul_res1[8117],mul_res1[8118],mul_res1[8119],mul_res1[8120],mul_res1[8121],mul_res1[8122],mul_res1[8123],mul_res1[8124],mul_res1[8125],mul_res1[8126],mul_res1[8127],mul_res1[8128],mul_res1[8129],mul_res1[8130],mul_res1[8131],mul_res1[8132],mul_res1[8133],mul_res1[8134],mul_res1[8135],mul_res1[8136],mul_res1[8137],mul_res1[8138],mul_res1[8139],mul_res1[8140],mul_res1[8141],mul_res1[8142],mul_res1[8143],mul_res1[8144],mul_res1[8145],mul_res1[8146],mul_res1[8147],mul_res1[8148],mul_res1[8149],mul_res1[8150],mul_res1[8151],mul_res1[8152],mul_res1[8153],mul_res1[8154],mul_res1[8155],mul_res1[8156],mul_res1[8157],mul_res1[8158],mul_res1[8159],mul_res1[8160],mul_res1[8161],mul_res1[8162],mul_res1[8163],mul_res1[8164],mul_res1[8165],mul_res1[8166],mul_res1[8167],mul_res1[8168],mul_res1[8169],mul_res1[8170],mul_res1[8171],mul_res1[8172],mul_res1[8173],mul_res1[8174],mul_res1[8175],mul_res1[8176],mul_res1[8177],mul_res1[8178],mul_res1[8179],mul_res1[8180],mul_res1[8181],mul_res1[8182],mul_res1[8183],mul_res1[8184],mul_res1[8185],mul_res1[8186],mul_res1[8187],mul_res1[8188],mul_res1[8189],mul_res1[8190],mul_res1[8191],mul_res1[8192],mul_res1[8193],mul_res1[8194],mul_res1[8195],mul_res1[8196],mul_res1[8197],mul_res1[8198],mul_res1[8199],result_fc1[40]);


adder_200in adder_200in_mod_41(clk,rst,mul_res1[8200],mul_res1[8201],mul_res1[8202],mul_res1[8203],mul_res1[8204],mul_res1[8205],mul_res1[8206],mul_res1[8207],mul_res1[8208],mul_res1[8209],mul_res1[8210],mul_res1[8211],mul_res1[8212],mul_res1[8213],mul_res1[8214],mul_res1[8215],mul_res1[8216],mul_res1[8217],mul_res1[8218],mul_res1[8219],mul_res1[8220],mul_res1[8221],mul_res1[8222],mul_res1[8223],mul_res1[8224],mul_res1[8225],mul_res1[8226],mul_res1[8227],mul_res1[8228],mul_res1[8229],mul_res1[8230],mul_res1[8231],mul_res1[8232],mul_res1[8233],mul_res1[8234],mul_res1[8235],mul_res1[8236],mul_res1[8237],mul_res1[8238],mul_res1[8239],mul_res1[8240],mul_res1[8241],mul_res1[8242],mul_res1[8243],mul_res1[8244],mul_res1[8245],mul_res1[8246],mul_res1[8247],mul_res1[8248],mul_res1[8249],mul_res1[8250],mul_res1[8251],mul_res1[8252],mul_res1[8253],mul_res1[8254],mul_res1[8255],mul_res1[8256],mul_res1[8257],mul_res1[8258],mul_res1[8259],mul_res1[8260],mul_res1[8261],mul_res1[8262],mul_res1[8263],mul_res1[8264],mul_res1[8265],mul_res1[8266],mul_res1[8267],mul_res1[8268],mul_res1[8269],mul_res1[8270],mul_res1[8271],mul_res1[8272],mul_res1[8273],mul_res1[8274],mul_res1[8275],mul_res1[8276],mul_res1[8277],mul_res1[8278],mul_res1[8279],mul_res1[8280],mul_res1[8281],mul_res1[8282],mul_res1[8283],mul_res1[8284],mul_res1[8285],mul_res1[8286],mul_res1[8287],mul_res1[8288],mul_res1[8289],mul_res1[8290],mul_res1[8291],mul_res1[8292],mul_res1[8293],mul_res1[8294],mul_res1[8295],mul_res1[8296],mul_res1[8297],mul_res1[8298],mul_res1[8299],mul_res1[8300],mul_res1[8301],mul_res1[8302],mul_res1[8303],mul_res1[8304],mul_res1[8305],mul_res1[8306],mul_res1[8307],mul_res1[8308],mul_res1[8309],mul_res1[8310],mul_res1[8311],mul_res1[8312],mul_res1[8313],mul_res1[8314],mul_res1[8315],mul_res1[8316],mul_res1[8317],mul_res1[8318],mul_res1[8319],mul_res1[8320],mul_res1[8321],mul_res1[8322],mul_res1[8323],mul_res1[8324],mul_res1[8325],mul_res1[8326],mul_res1[8327],mul_res1[8328],mul_res1[8329],mul_res1[8330],mul_res1[8331],mul_res1[8332],mul_res1[8333],mul_res1[8334],mul_res1[8335],mul_res1[8336],mul_res1[8337],mul_res1[8338],mul_res1[8339],mul_res1[8340],mul_res1[8341],mul_res1[8342],mul_res1[8343],mul_res1[8344],mul_res1[8345],mul_res1[8346],mul_res1[8347],mul_res1[8348],mul_res1[8349],mul_res1[8350],mul_res1[8351],mul_res1[8352],mul_res1[8353],mul_res1[8354],mul_res1[8355],mul_res1[8356],mul_res1[8357],mul_res1[8358],mul_res1[8359],mul_res1[8360],mul_res1[8361],mul_res1[8362],mul_res1[8363],mul_res1[8364],mul_res1[8365],mul_res1[8366],mul_res1[8367],mul_res1[8368],mul_res1[8369],mul_res1[8370],mul_res1[8371],mul_res1[8372],mul_res1[8373],mul_res1[8374],mul_res1[8375],mul_res1[8376],mul_res1[8377],mul_res1[8378],mul_res1[8379],mul_res1[8380],mul_res1[8381],mul_res1[8382],mul_res1[8383],mul_res1[8384],mul_res1[8385],mul_res1[8386],mul_res1[8387],mul_res1[8388],mul_res1[8389],mul_res1[8390],mul_res1[8391],mul_res1[8392],mul_res1[8393],mul_res1[8394],mul_res1[8395],mul_res1[8396],mul_res1[8397],mul_res1[8398],mul_res1[8399],result_fc1[41]);


adder_200in adder_200in_mod_42(clk,rst,mul_res1[8400],mul_res1[8401],mul_res1[8402],mul_res1[8403],mul_res1[8404],mul_res1[8405],mul_res1[8406],mul_res1[8407],mul_res1[8408],mul_res1[8409],mul_res1[8410],mul_res1[8411],mul_res1[8412],mul_res1[8413],mul_res1[8414],mul_res1[8415],mul_res1[8416],mul_res1[8417],mul_res1[8418],mul_res1[8419],mul_res1[8420],mul_res1[8421],mul_res1[8422],mul_res1[8423],mul_res1[8424],mul_res1[8425],mul_res1[8426],mul_res1[8427],mul_res1[8428],mul_res1[8429],mul_res1[8430],mul_res1[8431],mul_res1[8432],mul_res1[8433],mul_res1[8434],mul_res1[8435],mul_res1[8436],mul_res1[8437],mul_res1[8438],mul_res1[8439],mul_res1[8440],mul_res1[8441],mul_res1[8442],mul_res1[8443],mul_res1[8444],mul_res1[8445],mul_res1[8446],mul_res1[8447],mul_res1[8448],mul_res1[8449],mul_res1[8450],mul_res1[8451],mul_res1[8452],mul_res1[8453],mul_res1[8454],mul_res1[8455],mul_res1[8456],mul_res1[8457],mul_res1[8458],mul_res1[8459],mul_res1[8460],mul_res1[8461],mul_res1[8462],mul_res1[8463],mul_res1[8464],mul_res1[8465],mul_res1[8466],mul_res1[8467],mul_res1[8468],mul_res1[8469],mul_res1[8470],mul_res1[8471],mul_res1[8472],mul_res1[8473],mul_res1[8474],mul_res1[8475],mul_res1[8476],mul_res1[8477],mul_res1[8478],mul_res1[8479],mul_res1[8480],mul_res1[8481],mul_res1[8482],mul_res1[8483],mul_res1[8484],mul_res1[8485],mul_res1[8486],mul_res1[8487],mul_res1[8488],mul_res1[8489],mul_res1[8490],mul_res1[8491],mul_res1[8492],mul_res1[8493],mul_res1[8494],mul_res1[8495],mul_res1[8496],mul_res1[8497],mul_res1[8498],mul_res1[8499],mul_res1[8500],mul_res1[8501],mul_res1[8502],mul_res1[8503],mul_res1[8504],mul_res1[8505],mul_res1[8506],mul_res1[8507],mul_res1[8508],mul_res1[8509],mul_res1[8510],mul_res1[8511],mul_res1[8512],mul_res1[8513],mul_res1[8514],mul_res1[8515],mul_res1[8516],mul_res1[8517],mul_res1[8518],mul_res1[8519],mul_res1[8520],mul_res1[8521],mul_res1[8522],mul_res1[8523],mul_res1[8524],mul_res1[8525],mul_res1[8526],mul_res1[8527],mul_res1[8528],mul_res1[8529],mul_res1[8530],mul_res1[8531],mul_res1[8532],mul_res1[8533],mul_res1[8534],mul_res1[8535],mul_res1[8536],mul_res1[8537],mul_res1[8538],mul_res1[8539],mul_res1[8540],mul_res1[8541],mul_res1[8542],mul_res1[8543],mul_res1[8544],mul_res1[8545],mul_res1[8546],mul_res1[8547],mul_res1[8548],mul_res1[8549],mul_res1[8550],mul_res1[8551],mul_res1[8552],mul_res1[8553],mul_res1[8554],mul_res1[8555],mul_res1[8556],mul_res1[8557],mul_res1[8558],mul_res1[8559],mul_res1[8560],mul_res1[8561],mul_res1[8562],mul_res1[8563],mul_res1[8564],mul_res1[8565],mul_res1[8566],mul_res1[8567],mul_res1[8568],mul_res1[8569],mul_res1[8570],mul_res1[8571],mul_res1[8572],mul_res1[8573],mul_res1[8574],mul_res1[8575],mul_res1[8576],mul_res1[8577],mul_res1[8578],mul_res1[8579],mul_res1[8580],mul_res1[8581],mul_res1[8582],mul_res1[8583],mul_res1[8584],mul_res1[8585],mul_res1[8586],mul_res1[8587],mul_res1[8588],mul_res1[8589],mul_res1[8590],mul_res1[8591],mul_res1[8592],mul_res1[8593],mul_res1[8594],mul_res1[8595],mul_res1[8596],mul_res1[8597],mul_res1[8598],mul_res1[8599],result_fc1[42]);


adder_200in adder_200in_mod_43(clk,rst,mul_res1[8600],mul_res1[8601],mul_res1[8602],mul_res1[8603],mul_res1[8604],mul_res1[8605],mul_res1[8606],mul_res1[8607],mul_res1[8608],mul_res1[8609],mul_res1[8610],mul_res1[8611],mul_res1[8612],mul_res1[8613],mul_res1[8614],mul_res1[8615],mul_res1[8616],mul_res1[8617],mul_res1[8618],mul_res1[8619],mul_res1[8620],mul_res1[8621],mul_res1[8622],mul_res1[8623],mul_res1[8624],mul_res1[8625],mul_res1[8626],mul_res1[8627],mul_res1[8628],mul_res1[8629],mul_res1[8630],mul_res1[8631],mul_res1[8632],mul_res1[8633],mul_res1[8634],mul_res1[8635],mul_res1[8636],mul_res1[8637],mul_res1[8638],mul_res1[8639],mul_res1[8640],mul_res1[8641],mul_res1[8642],mul_res1[8643],mul_res1[8644],mul_res1[8645],mul_res1[8646],mul_res1[8647],mul_res1[8648],mul_res1[8649],mul_res1[8650],mul_res1[8651],mul_res1[8652],mul_res1[8653],mul_res1[8654],mul_res1[8655],mul_res1[8656],mul_res1[8657],mul_res1[8658],mul_res1[8659],mul_res1[8660],mul_res1[8661],mul_res1[8662],mul_res1[8663],mul_res1[8664],mul_res1[8665],mul_res1[8666],mul_res1[8667],mul_res1[8668],mul_res1[8669],mul_res1[8670],mul_res1[8671],mul_res1[8672],mul_res1[8673],mul_res1[8674],mul_res1[8675],mul_res1[8676],mul_res1[8677],mul_res1[8678],mul_res1[8679],mul_res1[8680],mul_res1[8681],mul_res1[8682],mul_res1[8683],mul_res1[8684],mul_res1[8685],mul_res1[8686],mul_res1[8687],mul_res1[8688],mul_res1[8689],mul_res1[8690],mul_res1[8691],mul_res1[8692],mul_res1[8693],mul_res1[8694],mul_res1[8695],mul_res1[8696],mul_res1[8697],mul_res1[8698],mul_res1[8699],mul_res1[8700],mul_res1[8701],mul_res1[8702],mul_res1[8703],mul_res1[8704],mul_res1[8705],mul_res1[8706],mul_res1[8707],mul_res1[8708],mul_res1[8709],mul_res1[8710],mul_res1[8711],mul_res1[8712],mul_res1[8713],mul_res1[8714],mul_res1[8715],mul_res1[8716],mul_res1[8717],mul_res1[8718],mul_res1[8719],mul_res1[8720],mul_res1[8721],mul_res1[8722],mul_res1[8723],mul_res1[8724],mul_res1[8725],mul_res1[8726],mul_res1[8727],mul_res1[8728],mul_res1[8729],mul_res1[8730],mul_res1[8731],mul_res1[8732],mul_res1[8733],mul_res1[8734],mul_res1[8735],mul_res1[8736],mul_res1[8737],mul_res1[8738],mul_res1[8739],mul_res1[8740],mul_res1[8741],mul_res1[8742],mul_res1[8743],mul_res1[8744],mul_res1[8745],mul_res1[8746],mul_res1[8747],mul_res1[8748],mul_res1[8749],mul_res1[8750],mul_res1[8751],mul_res1[8752],mul_res1[8753],mul_res1[8754],mul_res1[8755],mul_res1[8756],mul_res1[8757],mul_res1[8758],mul_res1[8759],mul_res1[8760],mul_res1[8761],mul_res1[8762],mul_res1[8763],mul_res1[8764],mul_res1[8765],mul_res1[8766],mul_res1[8767],mul_res1[8768],mul_res1[8769],mul_res1[8770],mul_res1[8771],mul_res1[8772],mul_res1[8773],mul_res1[8774],mul_res1[8775],mul_res1[8776],mul_res1[8777],mul_res1[8778],mul_res1[8779],mul_res1[8780],mul_res1[8781],mul_res1[8782],mul_res1[8783],mul_res1[8784],mul_res1[8785],mul_res1[8786],mul_res1[8787],mul_res1[8788],mul_res1[8789],mul_res1[8790],mul_res1[8791],mul_res1[8792],mul_res1[8793],mul_res1[8794],mul_res1[8795],mul_res1[8796],mul_res1[8797],mul_res1[8798],mul_res1[8799],result_fc1[43]);


adder_200in adder_200in_mod_44(clk,rst,mul_res1[8800],mul_res1[8801],mul_res1[8802],mul_res1[8803],mul_res1[8804],mul_res1[8805],mul_res1[8806],mul_res1[8807],mul_res1[8808],mul_res1[8809],mul_res1[8810],mul_res1[8811],mul_res1[8812],mul_res1[8813],mul_res1[8814],mul_res1[8815],mul_res1[8816],mul_res1[8817],mul_res1[8818],mul_res1[8819],mul_res1[8820],mul_res1[8821],mul_res1[8822],mul_res1[8823],mul_res1[8824],mul_res1[8825],mul_res1[8826],mul_res1[8827],mul_res1[8828],mul_res1[8829],mul_res1[8830],mul_res1[8831],mul_res1[8832],mul_res1[8833],mul_res1[8834],mul_res1[8835],mul_res1[8836],mul_res1[8837],mul_res1[8838],mul_res1[8839],mul_res1[8840],mul_res1[8841],mul_res1[8842],mul_res1[8843],mul_res1[8844],mul_res1[8845],mul_res1[8846],mul_res1[8847],mul_res1[8848],mul_res1[8849],mul_res1[8850],mul_res1[8851],mul_res1[8852],mul_res1[8853],mul_res1[8854],mul_res1[8855],mul_res1[8856],mul_res1[8857],mul_res1[8858],mul_res1[8859],mul_res1[8860],mul_res1[8861],mul_res1[8862],mul_res1[8863],mul_res1[8864],mul_res1[8865],mul_res1[8866],mul_res1[8867],mul_res1[8868],mul_res1[8869],mul_res1[8870],mul_res1[8871],mul_res1[8872],mul_res1[8873],mul_res1[8874],mul_res1[8875],mul_res1[8876],mul_res1[8877],mul_res1[8878],mul_res1[8879],mul_res1[8880],mul_res1[8881],mul_res1[8882],mul_res1[8883],mul_res1[8884],mul_res1[8885],mul_res1[8886],mul_res1[8887],mul_res1[8888],mul_res1[8889],mul_res1[8890],mul_res1[8891],mul_res1[8892],mul_res1[8893],mul_res1[8894],mul_res1[8895],mul_res1[8896],mul_res1[8897],mul_res1[8898],mul_res1[8899],mul_res1[8900],mul_res1[8901],mul_res1[8902],mul_res1[8903],mul_res1[8904],mul_res1[8905],mul_res1[8906],mul_res1[8907],mul_res1[8908],mul_res1[8909],mul_res1[8910],mul_res1[8911],mul_res1[8912],mul_res1[8913],mul_res1[8914],mul_res1[8915],mul_res1[8916],mul_res1[8917],mul_res1[8918],mul_res1[8919],mul_res1[8920],mul_res1[8921],mul_res1[8922],mul_res1[8923],mul_res1[8924],mul_res1[8925],mul_res1[8926],mul_res1[8927],mul_res1[8928],mul_res1[8929],mul_res1[8930],mul_res1[8931],mul_res1[8932],mul_res1[8933],mul_res1[8934],mul_res1[8935],mul_res1[8936],mul_res1[8937],mul_res1[8938],mul_res1[8939],mul_res1[8940],mul_res1[8941],mul_res1[8942],mul_res1[8943],mul_res1[8944],mul_res1[8945],mul_res1[8946],mul_res1[8947],mul_res1[8948],mul_res1[8949],mul_res1[8950],mul_res1[8951],mul_res1[8952],mul_res1[8953],mul_res1[8954],mul_res1[8955],mul_res1[8956],mul_res1[8957],mul_res1[8958],mul_res1[8959],mul_res1[8960],mul_res1[8961],mul_res1[8962],mul_res1[8963],mul_res1[8964],mul_res1[8965],mul_res1[8966],mul_res1[8967],mul_res1[8968],mul_res1[8969],mul_res1[8970],mul_res1[8971],mul_res1[8972],mul_res1[8973],mul_res1[8974],mul_res1[8975],mul_res1[8976],mul_res1[8977],mul_res1[8978],mul_res1[8979],mul_res1[8980],mul_res1[8981],mul_res1[8982],mul_res1[8983],mul_res1[8984],mul_res1[8985],mul_res1[8986],mul_res1[8987],mul_res1[8988],mul_res1[8989],mul_res1[8990],mul_res1[8991],mul_res1[8992],mul_res1[8993],mul_res1[8994],mul_res1[8995],mul_res1[8996],mul_res1[8997],mul_res1[8998],mul_res1[8999],result_fc1[44]);


adder_200in adder_200in_mod_45(clk,rst,mul_res1[9000],mul_res1[9001],mul_res1[9002],mul_res1[9003],mul_res1[9004],mul_res1[9005],mul_res1[9006],mul_res1[9007],mul_res1[9008],mul_res1[9009],mul_res1[9010],mul_res1[9011],mul_res1[9012],mul_res1[9013],mul_res1[9014],mul_res1[9015],mul_res1[9016],mul_res1[9017],mul_res1[9018],mul_res1[9019],mul_res1[9020],mul_res1[9021],mul_res1[9022],mul_res1[9023],mul_res1[9024],mul_res1[9025],mul_res1[9026],mul_res1[9027],mul_res1[9028],mul_res1[9029],mul_res1[9030],mul_res1[9031],mul_res1[9032],mul_res1[9033],mul_res1[9034],mul_res1[9035],mul_res1[9036],mul_res1[9037],mul_res1[9038],mul_res1[9039],mul_res1[9040],mul_res1[9041],mul_res1[9042],mul_res1[9043],mul_res1[9044],mul_res1[9045],mul_res1[9046],mul_res1[9047],mul_res1[9048],mul_res1[9049],mul_res1[9050],mul_res1[9051],mul_res1[9052],mul_res1[9053],mul_res1[9054],mul_res1[9055],mul_res1[9056],mul_res1[9057],mul_res1[9058],mul_res1[9059],mul_res1[9060],mul_res1[9061],mul_res1[9062],mul_res1[9063],mul_res1[9064],mul_res1[9065],mul_res1[9066],mul_res1[9067],mul_res1[9068],mul_res1[9069],mul_res1[9070],mul_res1[9071],mul_res1[9072],mul_res1[9073],mul_res1[9074],mul_res1[9075],mul_res1[9076],mul_res1[9077],mul_res1[9078],mul_res1[9079],mul_res1[9080],mul_res1[9081],mul_res1[9082],mul_res1[9083],mul_res1[9084],mul_res1[9085],mul_res1[9086],mul_res1[9087],mul_res1[9088],mul_res1[9089],mul_res1[9090],mul_res1[9091],mul_res1[9092],mul_res1[9093],mul_res1[9094],mul_res1[9095],mul_res1[9096],mul_res1[9097],mul_res1[9098],mul_res1[9099],mul_res1[9100],mul_res1[9101],mul_res1[9102],mul_res1[9103],mul_res1[9104],mul_res1[9105],mul_res1[9106],mul_res1[9107],mul_res1[9108],mul_res1[9109],mul_res1[9110],mul_res1[9111],mul_res1[9112],mul_res1[9113],mul_res1[9114],mul_res1[9115],mul_res1[9116],mul_res1[9117],mul_res1[9118],mul_res1[9119],mul_res1[9120],mul_res1[9121],mul_res1[9122],mul_res1[9123],mul_res1[9124],mul_res1[9125],mul_res1[9126],mul_res1[9127],mul_res1[9128],mul_res1[9129],mul_res1[9130],mul_res1[9131],mul_res1[9132],mul_res1[9133],mul_res1[9134],mul_res1[9135],mul_res1[9136],mul_res1[9137],mul_res1[9138],mul_res1[9139],mul_res1[9140],mul_res1[9141],mul_res1[9142],mul_res1[9143],mul_res1[9144],mul_res1[9145],mul_res1[9146],mul_res1[9147],mul_res1[9148],mul_res1[9149],mul_res1[9150],mul_res1[9151],mul_res1[9152],mul_res1[9153],mul_res1[9154],mul_res1[9155],mul_res1[9156],mul_res1[9157],mul_res1[9158],mul_res1[9159],mul_res1[9160],mul_res1[9161],mul_res1[9162],mul_res1[9163],mul_res1[9164],mul_res1[9165],mul_res1[9166],mul_res1[9167],mul_res1[9168],mul_res1[9169],mul_res1[9170],mul_res1[9171],mul_res1[9172],mul_res1[9173],mul_res1[9174],mul_res1[9175],mul_res1[9176],mul_res1[9177],mul_res1[9178],mul_res1[9179],mul_res1[9180],mul_res1[9181],mul_res1[9182],mul_res1[9183],mul_res1[9184],mul_res1[9185],mul_res1[9186],mul_res1[9187],mul_res1[9188],mul_res1[9189],mul_res1[9190],mul_res1[9191],mul_res1[9192],mul_res1[9193],mul_res1[9194],mul_res1[9195],mul_res1[9196],mul_res1[9197],mul_res1[9198],mul_res1[9199],result_fc1[45]);


adder_200in adder_200in_mod_46(clk,rst,mul_res1[9200],mul_res1[9201],mul_res1[9202],mul_res1[9203],mul_res1[9204],mul_res1[9205],mul_res1[9206],mul_res1[9207],mul_res1[9208],mul_res1[9209],mul_res1[9210],mul_res1[9211],mul_res1[9212],mul_res1[9213],mul_res1[9214],mul_res1[9215],mul_res1[9216],mul_res1[9217],mul_res1[9218],mul_res1[9219],mul_res1[9220],mul_res1[9221],mul_res1[9222],mul_res1[9223],mul_res1[9224],mul_res1[9225],mul_res1[9226],mul_res1[9227],mul_res1[9228],mul_res1[9229],mul_res1[9230],mul_res1[9231],mul_res1[9232],mul_res1[9233],mul_res1[9234],mul_res1[9235],mul_res1[9236],mul_res1[9237],mul_res1[9238],mul_res1[9239],mul_res1[9240],mul_res1[9241],mul_res1[9242],mul_res1[9243],mul_res1[9244],mul_res1[9245],mul_res1[9246],mul_res1[9247],mul_res1[9248],mul_res1[9249],mul_res1[9250],mul_res1[9251],mul_res1[9252],mul_res1[9253],mul_res1[9254],mul_res1[9255],mul_res1[9256],mul_res1[9257],mul_res1[9258],mul_res1[9259],mul_res1[9260],mul_res1[9261],mul_res1[9262],mul_res1[9263],mul_res1[9264],mul_res1[9265],mul_res1[9266],mul_res1[9267],mul_res1[9268],mul_res1[9269],mul_res1[9270],mul_res1[9271],mul_res1[9272],mul_res1[9273],mul_res1[9274],mul_res1[9275],mul_res1[9276],mul_res1[9277],mul_res1[9278],mul_res1[9279],mul_res1[9280],mul_res1[9281],mul_res1[9282],mul_res1[9283],mul_res1[9284],mul_res1[9285],mul_res1[9286],mul_res1[9287],mul_res1[9288],mul_res1[9289],mul_res1[9290],mul_res1[9291],mul_res1[9292],mul_res1[9293],mul_res1[9294],mul_res1[9295],mul_res1[9296],mul_res1[9297],mul_res1[9298],mul_res1[9299],mul_res1[9300],mul_res1[9301],mul_res1[9302],mul_res1[9303],mul_res1[9304],mul_res1[9305],mul_res1[9306],mul_res1[9307],mul_res1[9308],mul_res1[9309],mul_res1[9310],mul_res1[9311],mul_res1[9312],mul_res1[9313],mul_res1[9314],mul_res1[9315],mul_res1[9316],mul_res1[9317],mul_res1[9318],mul_res1[9319],mul_res1[9320],mul_res1[9321],mul_res1[9322],mul_res1[9323],mul_res1[9324],mul_res1[9325],mul_res1[9326],mul_res1[9327],mul_res1[9328],mul_res1[9329],mul_res1[9330],mul_res1[9331],mul_res1[9332],mul_res1[9333],mul_res1[9334],mul_res1[9335],mul_res1[9336],mul_res1[9337],mul_res1[9338],mul_res1[9339],mul_res1[9340],mul_res1[9341],mul_res1[9342],mul_res1[9343],mul_res1[9344],mul_res1[9345],mul_res1[9346],mul_res1[9347],mul_res1[9348],mul_res1[9349],mul_res1[9350],mul_res1[9351],mul_res1[9352],mul_res1[9353],mul_res1[9354],mul_res1[9355],mul_res1[9356],mul_res1[9357],mul_res1[9358],mul_res1[9359],mul_res1[9360],mul_res1[9361],mul_res1[9362],mul_res1[9363],mul_res1[9364],mul_res1[9365],mul_res1[9366],mul_res1[9367],mul_res1[9368],mul_res1[9369],mul_res1[9370],mul_res1[9371],mul_res1[9372],mul_res1[9373],mul_res1[9374],mul_res1[9375],mul_res1[9376],mul_res1[9377],mul_res1[9378],mul_res1[9379],mul_res1[9380],mul_res1[9381],mul_res1[9382],mul_res1[9383],mul_res1[9384],mul_res1[9385],mul_res1[9386],mul_res1[9387],mul_res1[9388],mul_res1[9389],mul_res1[9390],mul_res1[9391],mul_res1[9392],mul_res1[9393],mul_res1[9394],mul_res1[9395],mul_res1[9396],mul_res1[9397],mul_res1[9398],mul_res1[9399],result_fc1[46]);


adder_200in adder_200in_mod_47(clk,rst,mul_res1[9400],mul_res1[9401],mul_res1[9402],mul_res1[9403],mul_res1[9404],mul_res1[9405],mul_res1[9406],mul_res1[9407],mul_res1[9408],mul_res1[9409],mul_res1[9410],mul_res1[9411],mul_res1[9412],mul_res1[9413],mul_res1[9414],mul_res1[9415],mul_res1[9416],mul_res1[9417],mul_res1[9418],mul_res1[9419],mul_res1[9420],mul_res1[9421],mul_res1[9422],mul_res1[9423],mul_res1[9424],mul_res1[9425],mul_res1[9426],mul_res1[9427],mul_res1[9428],mul_res1[9429],mul_res1[9430],mul_res1[9431],mul_res1[9432],mul_res1[9433],mul_res1[9434],mul_res1[9435],mul_res1[9436],mul_res1[9437],mul_res1[9438],mul_res1[9439],mul_res1[9440],mul_res1[9441],mul_res1[9442],mul_res1[9443],mul_res1[9444],mul_res1[9445],mul_res1[9446],mul_res1[9447],mul_res1[9448],mul_res1[9449],mul_res1[9450],mul_res1[9451],mul_res1[9452],mul_res1[9453],mul_res1[9454],mul_res1[9455],mul_res1[9456],mul_res1[9457],mul_res1[9458],mul_res1[9459],mul_res1[9460],mul_res1[9461],mul_res1[9462],mul_res1[9463],mul_res1[9464],mul_res1[9465],mul_res1[9466],mul_res1[9467],mul_res1[9468],mul_res1[9469],mul_res1[9470],mul_res1[9471],mul_res1[9472],mul_res1[9473],mul_res1[9474],mul_res1[9475],mul_res1[9476],mul_res1[9477],mul_res1[9478],mul_res1[9479],mul_res1[9480],mul_res1[9481],mul_res1[9482],mul_res1[9483],mul_res1[9484],mul_res1[9485],mul_res1[9486],mul_res1[9487],mul_res1[9488],mul_res1[9489],mul_res1[9490],mul_res1[9491],mul_res1[9492],mul_res1[9493],mul_res1[9494],mul_res1[9495],mul_res1[9496],mul_res1[9497],mul_res1[9498],mul_res1[9499],mul_res1[9500],mul_res1[9501],mul_res1[9502],mul_res1[9503],mul_res1[9504],mul_res1[9505],mul_res1[9506],mul_res1[9507],mul_res1[9508],mul_res1[9509],mul_res1[9510],mul_res1[9511],mul_res1[9512],mul_res1[9513],mul_res1[9514],mul_res1[9515],mul_res1[9516],mul_res1[9517],mul_res1[9518],mul_res1[9519],mul_res1[9520],mul_res1[9521],mul_res1[9522],mul_res1[9523],mul_res1[9524],mul_res1[9525],mul_res1[9526],mul_res1[9527],mul_res1[9528],mul_res1[9529],mul_res1[9530],mul_res1[9531],mul_res1[9532],mul_res1[9533],mul_res1[9534],mul_res1[9535],mul_res1[9536],mul_res1[9537],mul_res1[9538],mul_res1[9539],mul_res1[9540],mul_res1[9541],mul_res1[9542],mul_res1[9543],mul_res1[9544],mul_res1[9545],mul_res1[9546],mul_res1[9547],mul_res1[9548],mul_res1[9549],mul_res1[9550],mul_res1[9551],mul_res1[9552],mul_res1[9553],mul_res1[9554],mul_res1[9555],mul_res1[9556],mul_res1[9557],mul_res1[9558],mul_res1[9559],mul_res1[9560],mul_res1[9561],mul_res1[9562],mul_res1[9563],mul_res1[9564],mul_res1[9565],mul_res1[9566],mul_res1[9567],mul_res1[9568],mul_res1[9569],mul_res1[9570],mul_res1[9571],mul_res1[9572],mul_res1[9573],mul_res1[9574],mul_res1[9575],mul_res1[9576],mul_res1[9577],mul_res1[9578],mul_res1[9579],mul_res1[9580],mul_res1[9581],mul_res1[9582],mul_res1[9583],mul_res1[9584],mul_res1[9585],mul_res1[9586],mul_res1[9587],mul_res1[9588],mul_res1[9589],mul_res1[9590],mul_res1[9591],mul_res1[9592],mul_res1[9593],mul_res1[9594],mul_res1[9595],mul_res1[9596],mul_res1[9597],mul_res1[9598],mul_res1[9599],result_fc1[47]);


adder_200in adder_200in_mod_48(clk,rst,mul_res1[9600],mul_res1[9601],mul_res1[9602],mul_res1[9603],mul_res1[9604],mul_res1[9605],mul_res1[9606],mul_res1[9607],mul_res1[9608],mul_res1[9609],mul_res1[9610],mul_res1[9611],mul_res1[9612],mul_res1[9613],mul_res1[9614],mul_res1[9615],mul_res1[9616],mul_res1[9617],mul_res1[9618],mul_res1[9619],mul_res1[9620],mul_res1[9621],mul_res1[9622],mul_res1[9623],mul_res1[9624],mul_res1[9625],mul_res1[9626],mul_res1[9627],mul_res1[9628],mul_res1[9629],mul_res1[9630],mul_res1[9631],mul_res1[9632],mul_res1[9633],mul_res1[9634],mul_res1[9635],mul_res1[9636],mul_res1[9637],mul_res1[9638],mul_res1[9639],mul_res1[9640],mul_res1[9641],mul_res1[9642],mul_res1[9643],mul_res1[9644],mul_res1[9645],mul_res1[9646],mul_res1[9647],mul_res1[9648],mul_res1[9649],mul_res1[9650],mul_res1[9651],mul_res1[9652],mul_res1[9653],mul_res1[9654],mul_res1[9655],mul_res1[9656],mul_res1[9657],mul_res1[9658],mul_res1[9659],mul_res1[9660],mul_res1[9661],mul_res1[9662],mul_res1[9663],mul_res1[9664],mul_res1[9665],mul_res1[9666],mul_res1[9667],mul_res1[9668],mul_res1[9669],mul_res1[9670],mul_res1[9671],mul_res1[9672],mul_res1[9673],mul_res1[9674],mul_res1[9675],mul_res1[9676],mul_res1[9677],mul_res1[9678],mul_res1[9679],mul_res1[9680],mul_res1[9681],mul_res1[9682],mul_res1[9683],mul_res1[9684],mul_res1[9685],mul_res1[9686],mul_res1[9687],mul_res1[9688],mul_res1[9689],mul_res1[9690],mul_res1[9691],mul_res1[9692],mul_res1[9693],mul_res1[9694],mul_res1[9695],mul_res1[9696],mul_res1[9697],mul_res1[9698],mul_res1[9699],mul_res1[9700],mul_res1[9701],mul_res1[9702],mul_res1[9703],mul_res1[9704],mul_res1[9705],mul_res1[9706],mul_res1[9707],mul_res1[9708],mul_res1[9709],mul_res1[9710],mul_res1[9711],mul_res1[9712],mul_res1[9713],mul_res1[9714],mul_res1[9715],mul_res1[9716],mul_res1[9717],mul_res1[9718],mul_res1[9719],mul_res1[9720],mul_res1[9721],mul_res1[9722],mul_res1[9723],mul_res1[9724],mul_res1[9725],mul_res1[9726],mul_res1[9727],mul_res1[9728],mul_res1[9729],mul_res1[9730],mul_res1[9731],mul_res1[9732],mul_res1[9733],mul_res1[9734],mul_res1[9735],mul_res1[9736],mul_res1[9737],mul_res1[9738],mul_res1[9739],mul_res1[9740],mul_res1[9741],mul_res1[9742],mul_res1[9743],mul_res1[9744],mul_res1[9745],mul_res1[9746],mul_res1[9747],mul_res1[9748],mul_res1[9749],mul_res1[9750],mul_res1[9751],mul_res1[9752],mul_res1[9753],mul_res1[9754],mul_res1[9755],mul_res1[9756],mul_res1[9757],mul_res1[9758],mul_res1[9759],mul_res1[9760],mul_res1[9761],mul_res1[9762],mul_res1[9763],mul_res1[9764],mul_res1[9765],mul_res1[9766],mul_res1[9767],mul_res1[9768],mul_res1[9769],mul_res1[9770],mul_res1[9771],mul_res1[9772],mul_res1[9773],mul_res1[9774],mul_res1[9775],mul_res1[9776],mul_res1[9777],mul_res1[9778],mul_res1[9779],mul_res1[9780],mul_res1[9781],mul_res1[9782],mul_res1[9783],mul_res1[9784],mul_res1[9785],mul_res1[9786],mul_res1[9787],mul_res1[9788],mul_res1[9789],mul_res1[9790],mul_res1[9791],mul_res1[9792],mul_res1[9793],mul_res1[9794],mul_res1[9795],mul_res1[9796],mul_res1[9797],mul_res1[9798],mul_res1[9799],result_fc1[48]);


adder_200in adder_200in_mod_49(clk,rst,mul_res1[9800],mul_res1[9801],mul_res1[9802],mul_res1[9803],mul_res1[9804],mul_res1[9805],mul_res1[9806],mul_res1[9807],mul_res1[9808],mul_res1[9809],mul_res1[9810],mul_res1[9811],mul_res1[9812],mul_res1[9813],mul_res1[9814],mul_res1[9815],mul_res1[9816],mul_res1[9817],mul_res1[9818],mul_res1[9819],mul_res1[9820],mul_res1[9821],mul_res1[9822],mul_res1[9823],mul_res1[9824],mul_res1[9825],mul_res1[9826],mul_res1[9827],mul_res1[9828],mul_res1[9829],mul_res1[9830],mul_res1[9831],mul_res1[9832],mul_res1[9833],mul_res1[9834],mul_res1[9835],mul_res1[9836],mul_res1[9837],mul_res1[9838],mul_res1[9839],mul_res1[9840],mul_res1[9841],mul_res1[9842],mul_res1[9843],mul_res1[9844],mul_res1[9845],mul_res1[9846],mul_res1[9847],mul_res1[9848],mul_res1[9849],mul_res1[9850],mul_res1[9851],mul_res1[9852],mul_res1[9853],mul_res1[9854],mul_res1[9855],mul_res1[9856],mul_res1[9857],mul_res1[9858],mul_res1[9859],mul_res1[9860],mul_res1[9861],mul_res1[9862],mul_res1[9863],mul_res1[9864],mul_res1[9865],mul_res1[9866],mul_res1[9867],mul_res1[9868],mul_res1[9869],mul_res1[9870],mul_res1[9871],mul_res1[9872],mul_res1[9873],mul_res1[9874],mul_res1[9875],mul_res1[9876],mul_res1[9877],mul_res1[9878],mul_res1[9879],mul_res1[9880],mul_res1[9881],mul_res1[9882],mul_res1[9883],mul_res1[9884],mul_res1[9885],mul_res1[9886],mul_res1[9887],mul_res1[9888],mul_res1[9889],mul_res1[9890],mul_res1[9891],mul_res1[9892],mul_res1[9893],mul_res1[9894],mul_res1[9895],mul_res1[9896],mul_res1[9897],mul_res1[9898],mul_res1[9899],mul_res1[9900],mul_res1[9901],mul_res1[9902],mul_res1[9903],mul_res1[9904],mul_res1[9905],mul_res1[9906],mul_res1[9907],mul_res1[9908],mul_res1[9909],mul_res1[9910],mul_res1[9911],mul_res1[9912],mul_res1[9913],mul_res1[9914],mul_res1[9915],mul_res1[9916],mul_res1[9917],mul_res1[9918],mul_res1[9919],mul_res1[9920],mul_res1[9921],mul_res1[9922],mul_res1[9923],mul_res1[9924],mul_res1[9925],mul_res1[9926],mul_res1[9927],mul_res1[9928],mul_res1[9929],mul_res1[9930],mul_res1[9931],mul_res1[9932],mul_res1[9933],mul_res1[9934],mul_res1[9935],mul_res1[9936],mul_res1[9937],mul_res1[9938],mul_res1[9939],mul_res1[9940],mul_res1[9941],mul_res1[9942],mul_res1[9943],mul_res1[9944],mul_res1[9945],mul_res1[9946],mul_res1[9947],mul_res1[9948],mul_res1[9949],mul_res1[9950],mul_res1[9951],mul_res1[9952],mul_res1[9953],mul_res1[9954],mul_res1[9955],mul_res1[9956],mul_res1[9957],mul_res1[9958],mul_res1[9959],mul_res1[9960],mul_res1[9961],mul_res1[9962],mul_res1[9963],mul_res1[9964],mul_res1[9965],mul_res1[9966],mul_res1[9967],mul_res1[9968],mul_res1[9969],mul_res1[9970],mul_res1[9971],mul_res1[9972],mul_res1[9973],mul_res1[9974],mul_res1[9975],mul_res1[9976],mul_res1[9977],mul_res1[9978],mul_res1[9979],mul_res1[9980],mul_res1[9981],mul_res1[9982],mul_res1[9983],mul_res1[9984],mul_res1[9985],mul_res1[9986],mul_res1[9987],mul_res1[9988],mul_res1[9989],mul_res1[9990],mul_res1[9991],mul_res1[9992],mul_res1[9993],mul_res1[9994],mul_res1[9995],mul_res1[9996],mul_res1[9997],mul_res1[9998],mul_res1[9999],result_fc1[49]);


adder_200in adder_200in_mod_50(clk,rst,mul_res1[10000],mul_res1[10001],mul_res1[10002],mul_res1[10003],mul_res1[10004],mul_res1[10005],mul_res1[10006],mul_res1[10007],mul_res1[10008],mul_res1[10009],mul_res1[10010],mul_res1[10011],mul_res1[10012],mul_res1[10013],mul_res1[10014],mul_res1[10015],mul_res1[10016],mul_res1[10017],mul_res1[10018],mul_res1[10019],mul_res1[10020],mul_res1[10021],mul_res1[10022],mul_res1[10023],mul_res1[10024],mul_res1[10025],mul_res1[10026],mul_res1[10027],mul_res1[10028],mul_res1[10029],mul_res1[10030],mul_res1[10031],mul_res1[10032],mul_res1[10033],mul_res1[10034],mul_res1[10035],mul_res1[10036],mul_res1[10037],mul_res1[10038],mul_res1[10039],mul_res1[10040],mul_res1[10041],mul_res1[10042],mul_res1[10043],mul_res1[10044],mul_res1[10045],mul_res1[10046],mul_res1[10047],mul_res1[10048],mul_res1[10049],mul_res1[10050],mul_res1[10051],mul_res1[10052],mul_res1[10053],mul_res1[10054],mul_res1[10055],mul_res1[10056],mul_res1[10057],mul_res1[10058],mul_res1[10059],mul_res1[10060],mul_res1[10061],mul_res1[10062],mul_res1[10063],mul_res1[10064],mul_res1[10065],mul_res1[10066],mul_res1[10067],mul_res1[10068],mul_res1[10069],mul_res1[10070],mul_res1[10071],mul_res1[10072],mul_res1[10073],mul_res1[10074],mul_res1[10075],mul_res1[10076],mul_res1[10077],mul_res1[10078],mul_res1[10079],mul_res1[10080],mul_res1[10081],mul_res1[10082],mul_res1[10083],mul_res1[10084],mul_res1[10085],mul_res1[10086],mul_res1[10087],mul_res1[10088],mul_res1[10089],mul_res1[10090],mul_res1[10091],mul_res1[10092],mul_res1[10093],mul_res1[10094],mul_res1[10095],mul_res1[10096],mul_res1[10097],mul_res1[10098],mul_res1[10099],mul_res1[10100],mul_res1[10101],mul_res1[10102],mul_res1[10103],mul_res1[10104],mul_res1[10105],mul_res1[10106],mul_res1[10107],mul_res1[10108],mul_res1[10109],mul_res1[10110],mul_res1[10111],mul_res1[10112],mul_res1[10113],mul_res1[10114],mul_res1[10115],mul_res1[10116],mul_res1[10117],mul_res1[10118],mul_res1[10119],mul_res1[10120],mul_res1[10121],mul_res1[10122],mul_res1[10123],mul_res1[10124],mul_res1[10125],mul_res1[10126],mul_res1[10127],mul_res1[10128],mul_res1[10129],mul_res1[10130],mul_res1[10131],mul_res1[10132],mul_res1[10133],mul_res1[10134],mul_res1[10135],mul_res1[10136],mul_res1[10137],mul_res1[10138],mul_res1[10139],mul_res1[10140],mul_res1[10141],mul_res1[10142],mul_res1[10143],mul_res1[10144],mul_res1[10145],mul_res1[10146],mul_res1[10147],mul_res1[10148],mul_res1[10149],mul_res1[10150],mul_res1[10151],mul_res1[10152],mul_res1[10153],mul_res1[10154],mul_res1[10155],mul_res1[10156],mul_res1[10157],mul_res1[10158],mul_res1[10159],mul_res1[10160],mul_res1[10161],mul_res1[10162],mul_res1[10163],mul_res1[10164],mul_res1[10165],mul_res1[10166],mul_res1[10167],mul_res1[10168],mul_res1[10169],mul_res1[10170],mul_res1[10171],mul_res1[10172],mul_res1[10173],mul_res1[10174],mul_res1[10175],mul_res1[10176],mul_res1[10177],mul_res1[10178],mul_res1[10179],mul_res1[10180],mul_res1[10181],mul_res1[10182],mul_res1[10183],mul_res1[10184],mul_res1[10185],mul_res1[10186],mul_res1[10187],mul_res1[10188],mul_res1[10189],mul_res1[10190],mul_res1[10191],mul_res1[10192],mul_res1[10193],mul_res1[10194],mul_res1[10195],mul_res1[10196],mul_res1[10197],mul_res1[10198],mul_res1[10199],result_fc1[50]);


adder_200in adder_200in_mod_51(clk,rst,mul_res1[10200],mul_res1[10201],mul_res1[10202],mul_res1[10203],mul_res1[10204],mul_res1[10205],mul_res1[10206],mul_res1[10207],mul_res1[10208],mul_res1[10209],mul_res1[10210],mul_res1[10211],mul_res1[10212],mul_res1[10213],mul_res1[10214],mul_res1[10215],mul_res1[10216],mul_res1[10217],mul_res1[10218],mul_res1[10219],mul_res1[10220],mul_res1[10221],mul_res1[10222],mul_res1[10223],mul_res1[10224],mul_res1[10225],mul_res1[10226],mul_res1[10227],mul_res1[10228],mul_res1[10229],mul_res1[10230],mul_res1[10231],mul_res1[10232],mul_res1[10233],mul_res1[10234],mul_res1[10235],mul_res1[10236],mul_res1[10237],mul_res1[10238],mul_res1[10239],mul_res1[10240],mul_res1[10241],mul_res1[10242],mul_res1[10243],mul_res1[10244],mul_res1[10245],mul_res1[10246],mul_res1[10247],mul_res1[10248],mul_res1[10249],mul_res1[10250],mul_res1[10251],mul_res1[10252],mul_res1[10253],mul_res1[10254],mul_res1[10255],mul_res1[10256],mul_res1[10257],mul_res1[10258],mul_res1[10259],mul_res1[10260],mul_res1[10261],mul_res1[10262],mul_res1[10263],mul_res1[10264],mul_res1[10265],mul_res1[10266],mul_res1[10267],mul_res1[10268],mul_res1[10269],mul_res1[10270],mul_res1[10271],mul_res1[10272],mul_res1[10273],mul_res1[10274],mul_res1[10275],mul_res1[10276],mul_res1[10277],mul_res1[10278],mul_res1[10279],mul_res1[10280],mul_res1[10281],mul_res1[10282],mul_res1[10283],mul_res1[10284],mul_res1[10285],mul_res1[10286],mul_res1[10287],mul_res1[10288],mul_res1[10289],mul_res1[10290],mul_res1[10291],mul_res1[10292],mul_res1[10293],mul_res1[10294],mul_res1[10295],mul_res1[10296],mul_res1[10297],mul_res1[10298],mul_res1[10299],mul_res1[10300],mul_res1[10301],mul_res1[10302],mul_res1[10303],mul_res1[10304],mul_res1[10305],mul_res1[10306],mul_res1[10307],mul_res1[10308],mul_res1[10309],mul_res1[10310],mul_res1[10311],mul_res1[10312],mul_res1[10313],mul_res1[10314],mul_res1[10315],mul_res1[10316],mul_res1[10317],mul_res1[10318],mul_res1[10319],mul_res1[10320],mul_res1[10321],mul_res1[10322],mul_res1[10323],mul_res1[10324],mul_res1[10325],mul_res1[10326],mul_res1[10327],mul_res1[10328],mul_res1[10329],mul_res1[10330],mul_res1[10331],mul_res1[10332],mul_res1[10333],mul_res1[10334],mul_res1[10335],mul_res1[10336],mul_res1[10337],mul_res1[10338],mul_res1[10339],mul_res1[10340],mul_res1[10341],mul_res1[10342],mul_res1[10343],mul_res1[10344],mul_res1[10345],mul_res1[10346],mul_res1[10347],mul_res1[10348],mul_res1[10349],mul_res1[10350],mul_res1[10351],mul_res1[10352],mul_res1[10353],mul_res1[10354],mul_res1[10355],mul_res1[10356],mul_res1[10357],mul_res1[10358],mul_res1[10359],mul_res1[10360],mul_res1[10361],mul_res1[10362],mul_res1[10363],mul_res1[10364],mul_res1[10365],mul_res1[10366],mul_res1[10367],mul_res1[10368],mul_res1[10369],mul_res1[10370],mul_res1[10371],mul_res1[10372],mul_res1[10373],mul_res1[10374],mul_res1[10375],mul_res1[10376],mul_res1[10377],mul_res1[10378],mul_res1[10379],mul_res1[10380],mul_res1[10381],mul_res1[10382],mul_res1[10383],mul_res1[10384],mul_res1[10385],mul_res1[10386],mul_res1[10387],mul_res1[10388],mul_res1[10389],mul_res1[10390],mul_res1[10391],mul_res1[10392],mul_res1[10393],mul_res1[10394],mul_res1[10395],mul_res1[10396],mul_res1[10397],mul_res1[10398],mul_res1[10399],result_fc1[51]);


adder_200in adder_200in_mod_52(clk,rst,mul_res1[10400],mul_res1[10401],mul_res1[10402],mul_res1[10403],mul_res1[10404],mul_res1[10405],mul_res1[10406],mul_res1[10407],mul_res1[10408],mul_res1[10409],mul_res1[10410],mul_res1[10411],mul_res1[10412],mul_res1[10413],mul_res1[10414],mul_res1[10415],mul_res1[10416],mul_res1[10417],mul_res1[10418],mul_res1[10419],mul_res1[10420],mul_res1[10421],mul_res1[10422],mul_res1[10423],mul_res1[10424],mul_res1[10425],mul_res1[10426],mul_res1[10427],mul_res1[10428],mul_res1[10429],mul_res1[10430],mul_res1[10431],mul_res1[10432],mul_res1[10433],mul_res1[10434],mul_res1[10435],mul_res1[10436],mul_res1[10437],mul_res1[10438],mul_res1[10439],mul_res1[10440],mul_res1[10441],mul_res1[10442],mul_res1[10443],mul_res1[10444],mul_res1[10445],mul_res1[10446],mul_res1[10447],mul_res1[10448],mul_res1[10449],mul_res1[10450],mul_res1[10451],mul_res1[10452],mul_res1[10453],mul_res1[10454],mul_res1[10455],mul_res1[10456],mul_res1[10457],mul_res1[10458],mul_res1[10459],mul_res1[10460],mul_res1[10461],mul_res1[10462],mul_res1[10463],mul_res1[10464],mul_res1[10465],mul_res1[10466],mul_res1[10467],mul_res1[10468],mul_res1[10469],mul_res1[10470],mul_res1[10471],mul_res1[10472],mul_res1[10473],mul_res1[10474],mul_res1[10475],mul_res1[10476],mul_res1[10477],mul_res1[10478],mul_res1[10479],mul_res1[10480],mul_res1[10481],mul_res1[10482],mul_res1[10483],mul_res1[10484],mul_res1[10485],mul_res1[10486],mul_res1[10487],mul_res1[10488],mul_res1[10489],mul_res1[10490],mul_res1[10491],mul_res1[10492],mul_res1[10493],mul_res1[10494],mul_res1[10495],mul_res1[10496],mul_res1[10497],mul_res1[10498],mul_res1[10499],mul_res1[10500],mul_res1[10501],mul_res1[10502],mul_res1[10503],mul_res1[10504],mul_res1[10505],mul_res1[10506],mul_res1[10507],mul_res1[10508],mul_res1[10509],mul_res1[10510],mul_res1[10511],mul_res1[10512],mul_res1[10513],mul_res1[10514],mul_res1[10515],mul_res1[10516],mul_res1[10517],mul_res1[10518],mul_res1[10519],mul_res1[10520],mul_res1[10521],mul_res1[10522],mul_res1[10523],mul_res1[10524],mul_res1[10525],mul_res1[10526],mul_res1[10527],mul_res1[10528],mul_res1[10529],mul_res1[10530],mul_res1[10531],mul_res1[10532],mul_res1[10533],mul_res1[10534],mul_res1[10535],mul_res1[10536],mul_res1[10537],mul_res1[10538],mul_res1[10539],mul_res1[10540],mul_res1[10541],mul_res1[10542],mul_res1[10543],mul_res1[10544],mul_res1[10545],mul_res1[10546],mul_res1[10547],mul_res1[10548],mul_res1[10549],mul_res1[10550],mul_res1[10551],mul_res1[10552],mul_res1[10553],mul_res1[10554],mul_res1[10555],mul_res1[10556],mul_res1[10557],mul_res1[10558],mul_res1[10559],mul_res1[10560],mul_res1[10561],mul_res1[10562],mul_res1[10563],mul_res1[10564],mul_res1[10565],mul_res1[10566],mul_res1[10567],mul_res1[10568],mul_res1[10569],mul_res1[10570],mul_res1[10571],mul_res1[10572],mul_res1[10573],mul_res1[10574],mul_res1[10575],mul_res1[10576],mul_res1[10577],mul_res1[10578],mul_res1[10579],mul_res1[10580],mul_res1[10581],mul_res1[10582],mul_res1[10583],mul_res1[10584],mul_res1[10585],mul_res1[10586],mul_res1[10587],mul_res1[10588],mul_res1[10589],mul_res1[10590],mul_res1[10591],mul_res1[10592],mul_res1[10593],mul_res1[10594],mul_res1[10595],mul_res1[10596],mul_res1[10597],mul_res1[10598],mul_res1[10599],result_fc1[52]);


adder_200in adder_200in_mod_53(clk,rst,mul_res1[10600],mul_res1[10601],mul_res1[10602],mul_res1[10603],mul_res1[10604],mul_res1[10605],mul_res1[10606],mul_res1[10607],mul_res1[10608],mul_res1[10609],mul_res1[10610],mul_res1[10611],mul_res1[10612],mul_res1[10613],mul_res1[10614],mul_res1[10615],mul_res1[10616],mul_res1[10617],mul_res1[10618],mul_res1[10619],mul_res1[10620],mul_res1[10621],mul_res1[10622],mul_res1[10623],mul_res1[10624],mul_res1[10625],mul_res1[10626],mul_res1[10627],mul_res1[10628],mul_res1[10629],mul_res1[10630],mul_res1[10631],mul_res1[10632],mul_res1[10633],mul_res1[10634],mul_res1[10635],mul_res1[10636],mul_res1[10637],mul_res1[10638],mul_res1[10639],mul_res1[10640],mul_res1[10641],mul_res1[10642],mul_res1[10643],mul_res1[10644],mul_res1[10645],mul_res1[10646],mul_res1[10647],mul_res1[10648],mul_res1[10649],mul_res1[10650],mul_res1[10651],mul_res1[10652],mul_res1[10653],mul_res1[10654],mul_res1[10655],mul_res1[10656],mul_res1[10657],mul_res1[10658],mul_res1[10659],mul_res1[10660],mul_res1[10661],mul_res1[10662],mul_res1[10663],mul_res1[10664],mul_res1[10665],mul_res1[10666],mul_res1[10667],mul_res1[10668],mul_res1[10669],mul_res1[10670],mul_res1[10671],mul_res1[10672],mul_res1[10673],mul_res1[10674],mul_res1[10675],mul_res1[10676],mul_res1[10677],mul_res1[10678],mul_res1[10679],mul_res1[10680],mul_res1[10681],mul_res1[10682],mul_res1[10683],mul_res1[10684],mul_res1[10685],mul_res1[10686],mul_res1[10687],mul_res1[10688],mul_res1[10689],mul_res1[10690],mul_res1[10691],mul_res1[10692],mul_res1[10693],mul_res1[10694],mul_res1[10695],mul_res1[10696],mul_res1[10697],mul_res1[10698],mul_res1[10699],mul_res1[10700],mul_res1[10701],mul_res1[10702],mul_res1[10703],mul_res1[10704],mul_res1[10705],mul_res1[10706],mul_res1[10707],mul_res1[10708],mul_res1[10709],mul_res1[10710],mul_res1[10711],mul_res1[10712],mul_res1[10713],mul_res1[10714],mul_res1[10715],mul_res1[10716],mul_res1[10717],mul_res1[10718],mul_res1[10719],mul_res1[10720],mul_res1[10721],mul_res1[10722],mul_res1[10723],mul_res1[10724],mul_res1[10725],mul_res1[10726],mul_res1[10727],mul_res1[10728],mul_res1[10729],mul_res1[10730],mul_res1[10731],mul_res1[10732],mul_res1[10733],mul_res1[10734],mul_res1[10735],mul_res1[10736],mul_res1[10737],mul_res1[10738],mul_res1[10739],mul_res1[10740],mul_res1[10741],mul_res1[10742],mul_res1[10743],mul_res1[10744],mul_res1[10745],mul_res1[10746],mul_res1[10747],mul_res1[10748],mul_res1[10749],mul_res1[10750],mul_res1[10751],mul_res1[10752],mul_res1[10753],mul_res1[10754],mul_res1[10755],mul_res1[10756],mul_res1[10757],mul_res1[10758],mul_res1[10759],mul_res1[10760],mul_res1[10761],mul_res1[10762],mul_res1[10763],mul_res1[10764],mul_res1[10765],mul_res1[10766],mul_res1[10767],mul_res1[10768],mul_res1[10769],mul_res1[10770],mul_res1[10771],mul_res1[10772],mul_res1[10773],mul_res1[10774],mul_res1[10775],mul_res1[10776],mul_res1[10777],mul_res1[10778],mul_res1[10779],mul_res1[10780],mul_res1[10781],mul_res1[10782],mul_res1[10783],mul_res1[10784],mul_res1[10785],mul_res1[10786],mul_res1[10787],mul_res1[10788],mul_res1[10789],mul_res1[10790],mul_res1[10791],mul_res1[10792],mul_res1[10793],mul_res1[10794],mul_res1[10795],mul_res1[10796],mul_res1[10797],mul_res1[10798],mul_res1[10799],result_fc1[53]);


adder_200in adder_200in_mod_54(clk,rst,mul_res1[10800],mul_res1[10801],mul_res1[10802],mul_res1[10803],mul_res1[10804],mul_res1[10805],mul_res1[10806],mul_res1[10807],mul_res1[10808],mul_res1[10809],mul_res1[10810],mul_res1[10811],mul_res1[10812],mul_res1[10813],mul_res1[10814],mul_res1[10815],mul_res1[10816],mul_res1[10817],mul_res1[10818],mul_res1[10819],mul_res1[10820],mul_res1[10821],mul_res1[10822],mul_res1[10823],mul_res1[10824],mul_res1[10825],mul_res1[10826],mul_res1[10827],mul_res1[10828],mul_res1[10829],mul_res1[10830],mul_res1[10831],mul_res1[10832],mul_res1[10833],mul_res1[10834],mul_res1[10835],mul_res1[10836],mul_res1[10837],mul_res1[10838],mul_res1[10839],mul_res1[10840],mul_res1[10841],mul_res1[10842],mul_res1[10843],mul_res1[10844],mul_res1[10845],mul_res1[10846],mul_res1[10847],mul_res1[10848],mul_res1[10849],mul_res1[10850],mul_res1[10851],mul_res1[10852],mul_res1[10853],mul_res1[10854],mul_res1[10855],mul_res1[10856],mul_res1[10857],mul_res1[10858],mul_res1[10859],mul_res1[10860],mul_res1[10861],mul_res1[10862],mul_res1[10863],mul_res1[10864],mul_res1[10865],mul_res1[10866],mul_res1[10867],mul_res1[10868],mul_res1[10869],mul_res1[10870],mul_res1[10871],mul_res1[10872],mul_res1[10873],mul_res1[10874],mul_res1[10875],mul_res1[10876],mul_res1[10877],mul_res1[10878],mul_res1[10879],mul_res1[10880],mul_res1[10881],mul_res1[10882],mul_res1[10883],mul_res1[10884],mul_res1[10885],mul_res1[10886],mul_res1[10887],mul_res1[10888],mul_res1[10889],mul_res1[10890],mul_res1[10891],mul_res1[10892],mul_res1[10893],mul_res1[10894],mul_res1[10895],mul_res1[10896],mul_res1[10897],mul_res1[10898],mul_res1[10899],mul_res1[10900],mul_res1[10901],mul_res1[10902],mul_res1[10903],mul_res1[10904],mul_res1[10905],mul_res1[10906],mul_res1[10907],mul_res1[10908],mul_res1[10909],mul_res1[10910],mul_res1[10911],mul_res1[10912],mul_res1[10913],mul_res1[10914],mul_res1[10915],mul_res1[10916],mul_res1[10917],mul_res1[10918],mul_res1[10919],mul_res1[10920],mul_res1[10921],mul_res1[10922],mul_res1[10923],mul_res1[10924],mul_res1[10925],mul_res1[10926],mul_res1[10927],mul_res1[10928],mul_res1[10929],mul_res1[10930],mul_res1[10931],mul_res1[10932],mul_res1[10933],mul_res1[10934],mul_res1[10935],mul_res1[10936],mul_res1[10937],mul_res1[10938],mul_res1[10939],mul_res1[10940],mul_res1[10941],mul_res1[10942],mul_res1[10943],mul_res1[10944],mul_res1[10945],mul_res1[10946],mul_res1[10947],mul_res1[10948],mul_res1[10949],mul_res1[10950],mul_res1[10951],mul_res1[10952],mul_res1[10953],mul_res1[10954],mul_res1[10955],mul_res1[10956],mul_res1[10957],mul_res1[10958],mul_res1[10959],mul_res1[10960],mul_res1[10961],mul_res1[10962],mul_res1[10963],mul_res1[10964],mul_res1[10965],mul_res1[10966],mul_res1[10967],mul_res1[10968],mul_res1[10969],mul_res1[10970],mul_res1[10971],mul_res1[10972],mul_res1[10973],mul_res1[10974],mul_res1[10975],mul_res1[10976],mul_res1[10977],mul_res1[10978],mul_res1[10979],mul_res1[10980],mul_res1[10981],mul_res1[10982],mul_res1[10983],mul_res1[10984],mul_res1[10985],mul_res1[10986],mul_res1[10987],mul_res1[10988],mul_res1[10989],mul_res1[10990],mul_res1[10991],mul_res1[10992],mul_res1[10993],mul_res1[10994],mul_res1[10995],mul_res1[10996],mul_res1[10997],mul_res1[10998],mul_res1[10999],result_fc1[54]);


adder_200in adder_200in_mod_55(clk,rst,mul_res1[11000],mul_res1[11001],mul_res1[11002],mul_res1[11003],mul_res1[11004],mul_res1[11005],mul_res1[11006],mul_res1[11007],mul_res1[11008],mul_res1[11009],mul_res1[11010],mul_res1[11011],mul_res1[11012],mul_res1[11013],mul_res1[11014],mul_res1[11015],mul_res1[11016],mul_res1[11017],mul_res1[11018],mul_res1[11019],mul_res1[11020],mul_res1[11021],mul_res1[11022],mul_res1[11023],mul_res1[11024],mul_res1[11025],mul_res1[11026],mul_res1[11027],mul_res1[11028],mul_res1[11029],mul_res1[11030],mul_res1[11031],mul_res1[11032],mul_res1[11033],mul_res1[11034],mul_res1[11035],mul_res1[11036],mul_res1[11037],mul_res1[11038],mul_res1[11039],mul_res1[11040],mul_res1[11041],mul_res1[11042],mul_res1[11043],mul_res1[11044],mul_res1[11045],mul_res1[11046],mul_res1[11047],mul_res1[11048],mul_res1[11049],mul_res1[11050],mul_res1[11051],mul_res1[11052],mul_res1[11053],mul_res1[11054],mul_res1[11055],mul_res1[11056],mul_res1[11057],mul_res1[11058],mul_res1[11059],mul_res1[11060],mul_res1[11061],mul_res1[11062],mul_res1[11063],mul_res1[11064],mul_res1[11065],mul_res1[11066],mul_res1[11067],mul_res1[11068],mul_res1[11069],mul_res1[11070],mul_res1[11071],mul_res1[11072],mul_res1[11073],mul_res1[11074],mul_res1[11075],mul_res1[11076],mul_res1[11077],mul_res1[11078],mul_res1[11079],mul_res1[11080],mul_res1[11081],mul_res1[11082],mul_res1[11083],mul_res1[11084],mul_res1[11085],mul_res1[11086],mul_res1[11087],mul_res1[11088],mul_res1[11089],mul_res1[11090],mul_res1[11091],mul_res1[11092],mul_res1[11093],mul_res1[11094],mul_res1[11095],mul_res1[11096],mul_res1[11097],mul_res1[11098],mul_res1[11099],mul_res1[11100],mul_res1[11101],mul_res1[11102],mul_res1[11103],mul_res1[11104],mul_res1[11105],mul_res1[11106],mul_res1[11107],mul_res1[11108],mul_res1[11109],mul_res1[11110],mul_res1[11111],mul_res1[11112],mul_res1[11113],mul_res1[11114],mul_res1[11115],mul_res1[11116],mul_res1[11117],mul_res1[11118],mul_res1[11119],mul_res1[11120],mul_res1[11121],mul_res1[11122],mul_res1[11123],mul_res1[11124],mul_res1[11125],mul_res1[11126],mul_res1[11127],mul_res1[11128],mul_res1[11129],mul_res1[11130],mul_res1[11131],mul_res1[11132],mul_res1[11133],mul_res1[11134],mul_res1[11135],mul_res1[11136],mul_res1[11137],mul_res1[11138],mul_res1[11139],mul_res1[11140],mul_res1[11141],mul_res1[11142],mul_res1[11143],mul_res1[11144],mul_res1[11145],mul_res1[11146],mul_res1[11147],mul_res1[11148],mul_res1[11149],mul_res1[11150],mul_res1[11151],mul_res1[11152],mul_res1[11153],mul_res1[11154],mul_res1[11155],mul_res1[11156],mul_res1[11157],mul_res1[11158],mul_res1[11159],mul_res1[11160],mul_res1[11161],mul_res1[11162],mul_res1[11163],mul_res1[11164],mul_res1[11165],mul_res1[11166],mul_res1[11167],mul_res1[11168],mul_res1[11169],mul_res1[11170],mul_res1[11171],mul_res1[11172],mul_res1[11173],mul_res1[11174],mul_res1[11175],mul_res1[11176],mul_res1[11177],mul_res1[11178],mul_res1[11179],mul_res1[11180],mul_res1[11181],mul_res1[11182],mul_res1[11183],mul_res1[11184],mul_res1[11185],mul_res1[11186],mul_res1[11187],mul_res1[11188],mul_res1[11189],mul_res1[11190],mul_res1[11191],mul_res1[11192],mul_res1[11193],mul_res1[11194],mul_res1[11195],mul_res1[11196],mul_res1[11197],mul_res1[11198],mul_res1[11199],result_fc1[55]);


adder_200in adder_200in_mod_56(clk,rst,mul_res1[11200],mul_res1[11201],mul_res1[11202],mul_res1[11203],mul_res1[11204],mul_res1[11205],mul_res1[11206],mul_res1[11207],mul_res1[11208],mul_res1[11209],mul_res1[11210],mul_res1[11211],mul_res1[11212],mul_res1[11213],mul_res1[11214],mul_res1[11215],mul_res1[11216],mul_res1[11217],mul_res1[11218],mul_res1[11219],mul_res1[11220],mul_res1[11221],mul_res1[11222],mul_res1[11223],mul_res1[11224],mul_res1[11225],mul_res1[11226],mul_res1[11227],mul_res1[11228],mul_res1[11229],mul_res1[11230],mul_res1[11231],mul_res1[11232],mul_res1[11233],mul_res1[11234],mul_res1[11235],mul_res1[11236],mul_res1[11237],mul_res1[11238],mul_res1[11239],mul_res1[11240],mul_res1[11241],mul_res1[11242],mul_res1[11243],mul_res1[11244],mul_res1[11245],mul_res1[11246],mul_res1[11247],mul_res1[11248],mul_res1[11249],mul_res1[11250],mul_res1[11251],mul_res1[11252],mul_res1[11253],mul_res1[11254],mul_res1[11255],mul_res1[11256],mul_res1[11257],mul_res1[11258],mul_res1[11259],mul_res1[11260],mul_res1[11261],mul_res1[11262],mul_res1[11263],mul_res1[11264],mul_res1[11265],mul_res1[11266],mul_res1[11267],mul_res1[11268],mul_res1[11269],mul_res1[11270],mul_res1[11271],mul_res1[11272],mul_res1[11273],mul_res1[11274],mul_res1[11275],mul_res1[11276],mul_res1[11277],mul_res1[11278],mul_res1[11279],mul_res1[11280],mul_res1[11281],mul_res1[11282],mul_res1[11283],mul_res1[11284],mul_res1[11285],mul_res1[11286],mul_res1[11287],mul_res1[11288],mul_res1[11289],mul_res1[11290],mul_res1[11291],mul_res1[11292],mul_res1[11293],mul_res1[11294],mul_res1[11295],mul_res1[11296],mul_res1[11297],mul_res1[11298],mul_res1[11299],mul_res1[11300],mul_res1[11301],mul_res1[11302],mul_res1[11303],mul_res1[11304],mul_res1[11305],mul_res1[11306],mul_res1[11307],mul_res1[11308],mul_res1[11309],mul_res1[11310],mul_res1[11311],mul_res1[11312],mul_res1[11313],mul_res1[11314],mul_res1[11315],mul_res1[11316],mul_res1[11317],mul_res1[11318],mul_res1[11319],mul_res1[11320],mul_res1[11321],mul_res1[11322],mul_res1[11323],mul_res1[11324],mul_res1[11325],mul_res1[11326],mul_res1[11327],mul_res1[11328],mul_res1[11329],mul_res1[11330],mul_res1[11331],mul_res1[11332],mul_res1[11333],mul_res1[11334],mul_res1[11335],mul_res1[11336],mul_res1[11337],mul_res1[11338],mul_res1[11339],mul_res1[11340],mul_res1[11341],mul_res1[11342],mul_res1[11343],mul_res1[11344],mul_res1[11345],mul_res1[11346],mul_res1[11347],mul_res1[11348],mul_res1[11349],mul_res1[11350],mul_res1[11351],mul_res1[11352],mul_res1[11353],mul_res1[11354],mul_res1[11355],mul_res1[11356],mul_res1[11357],mul_res1[11358],mul_res1[11359],mul_res1[11360],mul_res1[11361],mul_res1[11362],mul_res1[11363],mul_res1[11364],mul_res1[11365],mul_res1[11366],mul_res1[11367],mul_res1[11368],mul_res1[11369],mul_res1[11370],mul_res1[11371],mul_res1[11372],mul_res1[11373],mul_res1[11374],mul_res1[11375],mul_res1[11376],mul_res1[11377],mul_res1[11378],mul_res1[11379],mul_res1[11380],mul_res1[11381],mul_res1[11382],mul_res1[11383],mul_res1[11384],mul_res1[11385],mul_res1[11386],mul_res1[11387],mul_res1[11388],mul_res1[11389],mul_res1[11390],mul_res1[11391],mul_res1[11392],mul_res1[11393],mul_res1[11394],mul_res1[11395],mul_res1[11396],mul_res1[11397],mul_res1[11398],mul_res1[11399],result_fc1[56]);


adder_200in adder_200in_mod_57(clk,rst,mul_res1[11400],mul_res1[11401],mul_res1[11402],mul_res1[11403],mul_res1[11404],mul_res1[11405],mul_res1[11406],mul_res1[11407],mul_res1[11408],mul_res1[11409],mul_res1[11410],mul_res1[11411],mul_res1[11412],mul_res1[11413],mul_res1[11414],mul_res1[11415],mul_res1[11416],mul_res1[11417],mul_res1[11418],mul_res1[11419],mul_res1[11420],mul_res1[11421],mul_res1[11422],mul_res1[11423],mul_res1[11424],mul_res1[11425],mul_res1[11426],mul_res1[11427],mul_res1[11428],mul_res1[11429],mul_res1[11430],mul_res1[11431],mul_res1[11432],mul_res1[11433],mul_res1[11434],mul_res1[11435],mul_res1[11436],mul_res1[11437],mul_res1[11438],mul_res1[11439],mul_res1[11440],mul_res1[11441],mul_res1[11442],mul_res1[11443],mul_res1[11444],mul_res1[11445],mul_res1[11446],mul_res1[11447],mul_res1[11448],mul_res1[11449],mul_res1[11450],mul_res1[11451],mul_res1[11452],mul_res1[11453],mul_res1[11454],mul_res1[11455],mul_res1[11456],mul_res1[11457],mul_res1[11458],mul_res1[11459],mul_res1[11460],mul_res1[11461],mul_res1[11462],mul_res1[11463],mul_res1[11464],mul_res1[11465],mul_res1[11466],mul_res1[11467],mul_res1[11468],mul_res1[11469],mul_res1[11470],mul_res1[11471],mul_res1[11472],mul_res1[11473],mul_res1[11474],mul_res1[11475],mul_res1[11476],mul_res1[11477],mul_res1[11478],mul_res1[11479],mul_res1[11480],mul_res1[11481],mul_res1[11482],mul_res1[11483],mul_res1[11484],mul_res1[11485],mul_res1[11486],mul_res1[11487],mul_res1[11488],mul_res1[11489],mul_res1[11490],mul_res1[11491],mul_res1[11492],mul_res1[11493],mul_res1[11494],mul_res1[11495],mul_res1[11496],mul_res1[11497],mul_res1[11498],mul_res1[11499],mul_res1[11500],mul_res1[11501],mul_res1[11502],mul_res1[11503],mul_res1[11504],mul_res1[11505],mul_res1[11506],mul_res1[11507],mul_res1[11508],mul_res1[11509],mul_res1[11510],mul_res1[11511],mul_res1[11512],mul_res1[11513],mul_res1[11514],mul_res1[11515],mul_res1[11516],mul_res1[11517],mul_res1[11518],mul_res1[11519],mul_res1[11520],mul_res1[11521],mul_res1[11522],mul_res1[11523],mul_res1[11524],mul_res1[11525],mul_res1[11526],mul_res1[11527],mul_res1[11528],mul_res1[11529],mul_res1[11530],mul_res1[11531],mul_res1[11532],mul_res1[11533],mul_res1[11534],mul_res1[11535],mul_res1[11536],mul_res1[11537],mul_res1[11538],mul_res1[11539],mul_res1[11540],mul_res1[11541],mul_res1[11542],mul_res1[11543],mul_res1[11544],mul_res1[11545],mul_res1[11546],mul_res1[11547],mul_res1[11548],mul_res1[11549],mul_res1[11550],mul_res1[11551],mul_res1[11552],mul_res1[11553],mul_res1[11554],mul_res1[11555],mul_res1[11556],mul_res1[11557],mul_res1[11558],mul_res1[11559],mul_res1[11560],mul_res1[11561],mul_res1[11562],mul_res1[11563],mul_res1[11564],mul_res1[11565],mul_res1[11566],mul_res1[11567],mul_res1[11568],mul_res1[11569],mul_res1[11570],mul_res1[11571],mul_res1[11572],mul_res1[11573],mul_res1[11574],mul_res1[11575],mul_res1[11576],mul_res1[11577],mul_res1[11578],mul_res1[11579],mul_res1[11580],mul_res1[11581],mul_res1[11582],mul_res1[11583],mul_res1[11584],mul_res1[11585],mul_res1[11586],mul_res1[11587],mul_res1[11588],mul_res1[11589],mul_res1[11590],mul_res1[11591],mul_res1[11592],mul_res1[11593],mul_res1[11594],mul_res1[11595],mul_res1[11596],mul_res1[11597],mul_res1[11598],mul_res1[11599],result_fc1[57]);


adder_200in adder_200in_mod_58(clk,rst,mul_res1[11600],mul_res1[11601],mul_res1[11602],mul_res1[11603],mul_res1[11604],mul_res1[11605],mul_res1[11606],mul_res1[11607],mul_res1[11608],mul_res1[11609],mul_res1[11610],mul_res1[11611],mul_res1[11612],mul_res1[11613],mul_res1[11614],mul_res1[11615],mul_res1[11616],mul_res1[11617],mul_res1[11618],mul_res1[11619],mul_res1[11620],mul_res1[11621],mul_res1[11622],mul_res1[11623],mul_res1[11624],mul_res1[11625],mul_res1[11626],mul_res1[11627],mul_res1[11628],mul_res1[11629],mul_res1[11630],mul_res1[11631],mul_res1[11632],mul_res1[11633],mul_res1[11634],mul_res1[11635],mul_res1[11636],mul_res1[11637],mul_res1[11638],mul_res1[11639],mul_res1[11640],mul_res1[11641],mul_res1[11642],mul_res1[11643],mul_res1[11644],mul_res1[11645],mul_res1[11646],mul_res1[11647],mul_res1[11648],mul_res1[11649],mul_res1[11650],mul_res1[11651],mul_res1[11652],mul_res1[11653],mul_res1[11654],mul_res1[11655],mul_res1[11656],mul_res1[11657],mul_res1[11658],mul_res1[11659],mul_res1[11660],mul_res1[11661],mul_res1[11662],mul_res1[11663],mul_res1[11664],mul_res1[11665],mul_res1[11666],mul_res1[11667],mul_res1[11668],mul_res1[11669],mul_res1[11670],mul_res1[11671],mul_res1[11672],mul_res1[11673],mul_res1[11674],mul_res1[11675],mul_res1[11676],mul_res1[11677],mul_res1[11678],mul_res1[11679],mul_res1[11680],mul_res1[11681],mul_res1[11682],mul_res1[11683],mul_res1[11684],mul_res1[11685],mul_res1[11686],mul_res1[11687],mul_res1[11688],mul_res1[11689],mul_res1[11690],mul_res1[11691],mul_res1[11692],mul_res1[11693],mul_res1[11694],mul_res1[11695],mul_res1[11696],mul_res1[11697],mul_res1[11698],mul_res1[11699],mul_res1[11700],mul_res1[11701],mul_res1[11702],mul_res1[11703],mul_res1[11704],mul_res1[11705],mul_res1[11706],mul_res1[11707],mul_res1[11708],mul_res1[11709],mul_res1[11710],mul_res1[11711],mul_res1[11712],mul_res1[11713],mul_res1[11714],mul_res1[11715],mul_res1[11716],mul_res1[11717],mul_res1[11718],mul_res1[11719],mul_res1[11720],mul_res1[11721],mul_res1[11722],mul_res1[11723],mul_res1[11724],mul_res1[11725],mul_res1[11726],mul_res1[11727],mul_res1[11728],mul_res1[11729],mul_res1[11730],mul_res1[11731],mul_res1[11732],mul_res1[11733],mul_res1[11734],mul_res1[11735],mul_res1[11736],mul_res1[11737],mul_res1[11738],mul_res1[11739],mul_res1[11740],mul_res1[11741],mul_res1[11742],mul_res1[11743],mul_res1[11744],mul_res1[11745],mul_res1[11746],mul_res1[11747],mul_res1[11748],mul_res1[11749],mul_res1[11750],mul_res1[11751],mul_res1[11752],mul_res1[11753],mul_res1[11754],mul_res1[11755],mul_res1[11756],mul_res1[11757],mul_res1[11758],mul_res1[11759],mul_res1[11760],mul_res1[11761],mul_res1[11762],mul_res1[11763],mul_res1[11764],mul_res1[11765],mul_res1[11766],mul_res1[11767],mul_res1[11768],mul_res1[11769],mul_res1[11770],mul_res1[11771],mul_res1[11772],mul_res1[11773],mul_res1[11774],mul_res1[11775],mul_res1[11776],mul_res1[11777],mul_res1[11778],mul_res1[11779],mul_res1[11780],mul_res1[11781],mul_res1[11782],mul_res1[11783],mul_res1[11784],mul_res1[11785],mul_res1[11786],mul_res1[11787],mul_res1[11788],mul_res1[11789],mul_res1[11790],mul_res1[11791],mul_res1[11792],mul_res1[11793],mul_res1[11794],mul_res1[11795],mul_res1[11796],mul_res1[11797],mul_res1[11798],mul_res1[11799],result_fc1[58]);


adder_200in adder_200in_mod_59(clk,rst,mul_res1[11800],mul_res1[11801],mul_res1[11802],mul_res1[11803],mul_res1[11804],mul_res1[11805],mul_res1[11806],mul_res1[11807],mul_res1[11808],mul_res1[11809],mul_res1[11810],mul_res1[11811],mul_res1[11812],mul_res1[11813],mul_res1[11814],mul_res1[11815],mul_res1[11816],mul_res1[11817],mul_res1[11818],mul_res1[11819],mul_res1[11820],mul_res1[11821],mul_res1[11822],mul_res1[11823],mul_res1[11824],mul_res1[11825],mul_res1[11826],mul_res1[11827],mul_res1[11828],mul_res1[11829],mul_res1[11830],mul_res1[11831],mul_res1[11832],mul_res1[11833],mul_res1[11834],mul_res1[11835],mul_res1[11836],mul_res1[11837],mul_res1[11838],mul_res1[11839],mul_res1[11840],mul_res1[11841],mul_res1[11842],mul_res1[11843],mul_res1[11844],mul_res1[11845],mul_res1[11846],mul_res1[11847],mul_res1[11848],mul_res1[11849],mul_res1[11850],mul_res1[11851],mul_res1[11852],mul_res1[11853],mul_res1[11854],mul_res1[11855],mul_res1[11856],mul_res1[11857],mul_res1[11858],mul_res1[11859],mul_res1[11860],mul_res1[11861],mul_res1[11862],mul_res1[11863],mul_res1[11864],mul_res1[11865],mul_res1[11866],mul_res1[11867],mul_res1[11868],mul_res1[11869],mul_res1[11870],mul_res1[11871],mul_res1[11872],mul_res1[11873],mul_res1[11874],mul_res1[11875],mul_res1[11876],mul_res1[11877],mul_res1[11878],mul_res1[11879],mul_res1[11880],mul_res1[11881],mul_res1[11882],mul_res1[11883],mul_res1[11884],mul_res1[11885],mul_res1[11886],mul_res1[11887],mul_res1[11888],mul_res1[11889],mul_res1[11890],mul_res1[11891],mul_res1[11892],mul_res1[11893],mul_res1[11894],mul_res1[11895],mul_res1[11896],mul_res1[11897],mul_res1[11898],mul_res1[11899],mul_res1[11900],mul_res1[11901],mul_res1[11902],mul_res1[11903],mul_res1[11904],mul_res1[11905],mul_res1[11906],mul_res1[11907],mul_res1[11908],mul_res1[11909],mul_res1[11910],mul_res1[11911],mul_res1[11912],mul_res1[11913],mul_res1[11914],mul_res1[11915],mul_res1[11916],mul_res1[11917],mul_res1[11918],mul_res1[11919],mul_res1[11920],mul_res1[11921],mul_res1[11922],mul_res1[11923],mul_res1[11924],mul_res1[11925],mul_res1[11926],mul_res1[11927],mul_res1[11928],mul_res1[11929],mul_res1[11930],mul_res1[11931],mul_res1[11932],mul_res1[11933],mul_res1[11934],mul_res1[11935],mul_res1[11936],mul_res1[11937],mul_res1[11938],mul_res1[11939],mul_res1[11940],mul_res1[11941],mul_res1[11942],mul_res1[11943],mul_res1[11944],mul_res1[11945],mul_res1[11946],mul_res1[11947],mul_res1[11948],mul_res1[11949],mul_res1[11950],mul_res1[11951],mul_res1[11952],mul_res1[11953],mul_res1[11954],mul_res1[11955],mul_res1[11956],mul_res1[11957],mul_res1[11958],mul_res1[11959],mul_res1[11960],mul_res1[11961],mul_res1[11962],mul_res1[11963],mul_res1[11964],mul_res1[11965],mul_res1[11966],mul_res1[11967],mul_res1[11968],mul_res1[11969],mul_res1[11970],mul_res1[11971],mul_res1[11972],mul_res1[11973],mul_res1[11974],mul_res1[11975],mul_res1[11976],mul_res1[11977],mul_res1[11978],mul_res1[11979],mul_res1[11980],mul_res1[11981],mul_res1[11982],mul_res1[11983],mul_res1[11984],mul_res1[11985],mul_res1[11986],mul_res1[11987],mul_res1[11988],mul_res1[11989],mul_res1[11990],mul_res1[11991],mul_res1[11992],mul_res1[11993],mul_res1[11994],mul_res1[11995],mul_res1[11996],mul_res1[11997],mul_res1[11998],mul_res1[11999],result_fc1[59]);


adder_200in adder_200in_mod_60(clk,rst,mul_res1[12000],mul_res1[12001],mul_res1[12002],mul_res1[12003],mul_res1[12004],mul_res1[12005],mul_res1[12006],mul_res1[12007],mul_res1[12008],mul_res1[12009],mul_res1[12010],mul_res1[12011],mul_res1[12012],mul_res1[12013],mul_res1[12014],mul_res1[12015],mul_res1[12016],mul_res1[12017],mul_res1[12018],mul_res1[12019],mul_res1[12020],mul_res1[12021],mul_res1[12022],mul_res1[12023],mul_res1[12024],mul_res1[12025],mul_res1[12026],mul_res1[12027],mul_res1[12028],mul_res1[12029],mul_res1[12030],mul_res1[12031],mul_res1[12032],mul_res1[12033],mul_res1[12034],mul_res1[12035],mul_res1[12036],mul_res1[12037],mul_res1[12038],mul_res1[12039],mul_res1[12040],mul_res1[12041],mul_res1[12042],mul_res1[12043],mul_res1[12044],mul_res1[12045],mul_res1[12046],mul_res1[12047],mul_res1[12048],mul_res1[12049],mul_res1[12050],mul_res1[12051],mul_res1[12052],mul_res1[12053],mul_res1[12054],mul_res1[12055],mul_res1[12056],mul_res1[12057],mul_res1[12058],mul_res1[12059],mul_res1[12060],mul_res1[12061],mul_res1[12062],mul_res1[12063],mul_res1[12064],mul_res1[12065],mul_res1[12066],mul_res1[12067],mul_res1[12068],mul_res1[12069],mul_res1[12070],mul_res1[12071],mul_res1[12072],mul_res1[12073],mul_res1[12074],mul_res1[12075],mul_res1[12076],mul_res1[12077],mul_res1[12078],mul_res1[12079],mul_res1[12080],mul_res1[12081],mul_res1[12082],mul_res1[12083],mul_res1[12084],mul_res1[12085],mul_res1[12086],mul_res1[12087],mul_res1[12088],mul_res1[12089],mul_res1[12090],mul_res1[12091],mul_res1[12092],mul_res1[12093],mul_res1[12094],mul_res1[12095],mul_res1[12096],mul_res1[12097],mul_res1[12098],mul_res1[12099],mul_res1[12100],mul_res1[12101],mul_res1[12102],mul_res1[12103],mul_res1[12104],mul_res1[12105],mul_res1[12106],mul_res1[12107],mul_res1[12108],mul_res1[12109],mul_res1[12110],mul_res1[12111],mul_res1[12112],mul_res1[12113],mul_res1[12114],mul_res1[12115],mul_res1[12116],mul_res1[12117],mul_res1[12118],mul_res1[12119],mul_res1[12120],mul_res1[12121],mul_res1[12122],mul_res1[12123],mul_res1[12124],mul_res1[12125],mul_res1[12126],mul_res1[12127],mul_res1[12128],mul_res1[12129],mul_res1[12130],mul_res1[12131],mul_res1[12132],mul_res1[12133],mul_res1[12134],mul_res1[12135],mul_res1[12136],mul_res1[12137],mul_res1[12138],mul_res1[12139],mul_res1[12140],mul_res1[12141],mul_res1[12142],mul_res1[12143],mul_res1[12144],mul_res1[12145],mul_res1[12146],mul_res1[12147],mul_res1[12148],mul_res1[12149],mul_res1[12150],mul_res1[12151],mul_res1[12152],mul_res1[12153],mul_res1[12154],mul_res1[12155],mul_res1[12156],mul_res1[12157],mul_res1[12158],mul_res1[12159],mul_res1[12160],mul_res1[12161],mul_res1[12162],mul_res1[12163],mul_res1[12164],mul_res1[12165],mul_res1[12166],mul_res1[12167],mul_res1[12168],mul_res1[12169],mul_res1[12170],mul_res1[12171],mul_res1[12172],mul_res1[12173],mul_res1[12174],mul_res1[12175],mul_res1[12176],mul_res1[12177],mul_res1[12178],mul_res1[12179],mul_res1[12180],mul_res1[12181],mul_res1[12182],mul_res1[12183],mul_res1[12184],mul_res1[12185],mul_res1[12186],mul_res1[12187],mul_res1[12188],mul_res1[12189],mul_res1[12190],mul_res1[12191],mul_res1[12192],mul_res1[12193],mul_res1[12194],mul_res1[12195],mul_res1[12196],mul_res1[12197],mul_res1[12198],mul_res1[12199],result_fc1[60]);


adder_200in adder_200in_mod_61(clk,rst,mul_res1[12200],mul_res1[12201],mul_res1[12202],mul_res1[12203],mul_res1[12204],mul_res1[12205],mul_res1[12206],mul_res1[12207],mul_res1[12208],mul_res1[12209],mul_res1[12210],mul_res1[12211],mul_res1[12212],mul_res1[12213],mul_res1[12214],mul_res1[12215],mul_res1[12216],mul_res1[12217],mul_res1[12218],mul_res1[12219],mul_res1[12220],mul_res1[12221],mul_res1[12222],mul_res1[12223],mul_res1[12224],mul_res1[12225],mul_res1[12226],mul_res1[12227],mul_res1[12228],mul_res1[12229],mul_res1[12230],mul_res1[12231],mul_res1[12232],mul_res1[12233],mul_res1[12234],mul_res1[12235],mul_res1[12236],mul_res1[12237],mul_res1[12238],mul_res1[12239],mul_res1[12240],mul_res1[12241],mul_res1[12242],mul_res1[12243],mul_res1[12244],mul_res1[12245],mul_res1[12246],mul_res1[12247],mul_res1[12248],mul_res1[12249],mul_res1[12250],mul_res1[12251],mul_res1[12252],mul_res1[12253],mul_res1[12254],mul_res1[12255],mul_res1[12256],mul_res1[12257],mul_res1[12258],mul_res1[12259],mul_res1[12260],mul_res1[12261],mul_res1[12262],mul_res1[12263],mul_res1[12264],mul_res1[12265],mul_res1[12266],mul_res1[12267],mul_res1[12268],mul_res1[12269],mul_res1[12270],mul_res1[12271],mul_res1[12272],mul_res1[12273],mul_res1[12274],mul_res1[12275],mul_res1[12276],mul_res1[12277],mul_res1[12278],mul_res1[12279],mul_res1[12280],mul_res1[12281],mul_res1[12282],mul_res1[12283],mul_res1[12284],mul_res1[12285],mul_res1[12286],mul_res1[12287],mul_res1[12288],mul_res1[12289],mul_res1[12290],mul_res1[12291],mul_res1[12292],mul_res1[12293],mul_res1[12294],mul_res1[12295],mul_res1[12296],mul_res1[12297],mul_res1[12298],mul_res1[12299],mul_res1[12300],mul_res1[12301],mul_res1[12302],mul_res1[12303],mul_res1[12304],mul_res1[12305],mul_res1[12306],mul_res1[12307],mul_res1[12308],mul_res1[12309],mul_res1[12310],mul_res1[12311],mul_res1[12312],mul_res1[12313],mul_res1[12314],mul_res1[12315],mul_res1[12316],mul_res1[12317],mul_res1[12318],mul_res1[12319],mul_res1[12320],mul_res1[12321],mul_res1[12322],mul_res1[12323],mul_res1[12324],mul_res1[12325],mul_res1[12326],mul_res1[12327],mul_res1[12328],mul_res1[12329],mul_res1[12330],mul_res1[12331],mul_res1[12332],mul_res1[12333],mul_res1[12334],mul_res1[12335],mul_res1[12336],mul_res1[12337],mul_res1[12338],mul_res1[12339],mul_res1[12340],mul_res1[12341],mul_res1[12342],mul_res1[12343],mul_res1[12344],mul_res1[12345],mul_res1[12346],mul_res1[12347],mul_res1[12348],mul_res1[12349],mul_res1[12350],mul_res1[12351],mul_res1[12352],mul_res1[12353],mul_res1[12354],mul_res1[12355],mul_res1[12356],mul_res1[12357],mul_res1[12358],mul_res1[12359],mul_res1[12360],mul_res1[12361],mul_res1[12362],mul_res1[12363],mul_res1[12364],mul_res1[12365],mul_res1[12366],mul_res1[12367],mul_res1[12368],mul_res1[12369],mul_res1[12370],mul_res1[12371],mul_res1[12372],mul_res1[12373],mul_res1[12374],mul_res1[12375],mul_res1[12376],mul_res1[12377],mul_res1[12378],mul_res1[12379],mul_res1[12380],mul_res1[12381],mul_res1[12382],mul_res1[12383],mul_res1[12384],mul_res1[12385],mul_res1[12386],mul_res1[12387],mul_res1[12388],mul_res1[12389],mul_res1[12390],mul_res1[12391],mul_res1[12392],mul_res1[12393],mul_res1[12394],mul_res1[12395],mul_res1[12396],mul_res1[12397],mul_res1[12398],mul_res1[12399],result_fc1[61]);


adder_200in adder_200in_mod_62(clk,rst,mul_res1[12400],mul_res1[12401],mul_res1[12402],mul_res1[12403],mul_res1[12404],mul_res1[12405],mul_res1[12406],mul_res1[12407],mul_res1[12408],mul_res1[12409],mul_res1[12410],mul_res1[12411],mul_res1[12412],mul_res1[12413],mul_res1[12414],mul_res1[12415],mul_res1[12416],mul_res1[12417],mul_res1[12418],mul_res1[12419],mul_res1[12420],mul_res1[12421],mul_res1[12422],mul_res1[12423],mul_res1[12424],mul_res1[12425],mul_res1[12426],mul_res1[12427],mul_res1[12428],mul_res1[12429],mul_res1[12430],mul_res1[12431],mul_res1[12432],mul_res1[12433],mul_res1[12434],mul_res1[12435],mul_res1[12436],mul_res1[12437],mul_res1[12438],mul_res1[12439],mul_res1[12440],mul_res1[12441],mul_res1[12442],mul_res1[12443],mul_res1[12444],mul_res1[12445],mul_res1[12446],mul_res1[12447],mul_res1[12448],mul_res1[12449],mul_res1[12450],mul_res1[12451],mul_res1[12452],mul_res1[12453],mul_res1[12454],mul_res1[12455],mul_res1[12456],mul_res1[12457],mul_res1[12458],mul_res1[12459],mul_res1[12460],mul_res1[12461],mul_res1[12462],mul_res1[12463],mul_res1[12464],mul_res1[12465],mul_res1[12466],mul_res1[12467],mul_res1[12468],mul_res1[12469],mul_res1[12470],mul_res1[12471],mul_res1[12472],mul_res1[12473],mul_res1[12474],mul_res1[12475],mul_res1[12476],mul_res1[12477],mul_res1[12478],mul_res1[12479],mul_res1[12480],mul_res1[12481],mul_res1[12482],mul_res1[12483],mul_res1[12484],mul_res1[12485],mul_res1[12486],mul_res1[12487],mul_res1[12488],mul_res1[12489],mul_res1[12490],mul_res1[12491],mul_res1[12492],mul_res1[12493],mul_res1[12494],mul_res1[12495],mul_res1[12496],mul_res1[12497],mul_res1[12498],mul_res1[12499],mul_res1[12500],mul_res1[12501],mul_res1[12502],mul_res1[12503],mul_res1[12504],mul_res1[12505],mul_res1[12506],mul_res1[12507],mul_res1[12508],mul_res1[12509],mul_res1[12510],mul_res1[12511],mul_res1[12512],mul_res1[12513],mul_res1[12514],mul_res1[12515],mul_res1[12516],mul_res1[12517],mul_res1[12518],mul_res1[12519],mul_res1[12520],mul_res1[12521],mul_res1[12522],mul_res1[12523],mul_res1[12524],mul_res1[12525],mul_res1[12526],mul_res1[12527],mul_res1[12528],mul_res1[12529],mul_res1[12530],mul_res1[12531],mul_res1[12532],mul_res1[12533],mul_res1[12534],mul_res1[12535],mul_res1[12536],mul_res1[12537],mul_res1[12538],mul_res1[12539],mul_res1[12540],mul_res1[12541],mul_res1[12542],mul_res1[12543],mul_res1[12544],mul_res1[12545],mul_res1[12546],mul_res1[12547],mul_res1[12548],mul_res1[12549],mul_res1[12550],mul_res1[12551],mul_res1[12552],mul_res1[12553],mul_res1[12554],mul_res1[12555],mul_res1[12556],mul_res1[12557],mul_res1[12558],mul_res1[12559],mul_res1[12560],mul_res1[12561],mul_res1[12562],mul_res1[12563],mul_res1[12564],mul_res1[12565],mul_res1[12566],mul_res1[12567],mul_res1[12568],mul_res1[12569],mul_res1[12570],mul_res1[12571],mul_res1[12572],mul_res1[12573],mul_res1[12574],mul_res1[12575],mul_res1[12576],mul_res1[12577],mul_res1[12578],mul_res1[12579],mul_res1[12580],mul_res1[12581],mul_res1[12582],mul_res1[12583],mul_res1[12584],mul_res1[12585],mul_res1[12586],mul_res1[12587],mul_res1[12588],mul_res1[12589],mul_res1[12590],mul_res1[12591],mul_res1[12592],mul_res1[12593],mul_res1[12594],mul_res1[12595],mul_res1[12596],mul_res1[12597],mul_res1[12598],mul_res1[12599],result_fc1[62]);


adder_200in adder_200in_mod_63(clk,rst,mul_res1[12600],mul_res1[12601],mul_res1[12602],mul_res1[12603],mul_res1[12604],mul_res1[12605],mul_res1[12606],mul_res1[12607],mul_res1[12608],mul_res1[12609],mul_res1[12610],mul_res1[12611],mul_res1[12612],mul_res1[12613],mul_res1[12614],mul_res1[12615],mul_res1[12616],mul_res1[12617],mul_res1[12618],mul_res1[12619],mul_res1[12620],mul_res1[12621],mul_res1[12622],mul_res1[12623],mul_res1[12624],mul_res1[12625],mul_res1[12626],mul_res1[12627],mul_res1[12628],mul_res1[12629],mul_res1[12630],mul_res1[12631],mul_res1[12632],mul_res1[12633],mul_res1[12634],mul_res1[12635],mul_res1[12636],mul_res1[12637],mul_res1[12638],mul_res1[12639],mul_res1[12640],mul_res1[12641],mul_res1[12642],mul_res1[12643],mul_res1[12644],mul_res1[12645],mul_res1[12646],mul_res1[12647],mul_res1[12648],mul_res1[12649],mul_res1[12650],mul_res1[12651],mul_res1[12652],mul_res1[12653],mul_res1[12654],mul_res1[12655],mul_res1[12656],mul_res1[12657],mul_res1[12658],mul_res1[12659],mul_res1[12660],mul_res1[12661],mul_res1[12662],mul_res1[12663],mul_res1[12664],mul_res1[12665],mul_res1[12666],mul_res1[12667],mul_res1[12668],mul_res1[12669],mul_res1[12670],mul_res1[12671],mul_res1[12672],mul_res1[12673],mul_res1[12674],mul_res1[12675],mul_res1[12676],mul_res1[12677],mul_res1[12678],mul_res1[12679],mul_res1[12680],mul_res1[12681],mul_res1[12682],mul_res1[12683],mul_res1[12684],mul_res1[12685],mul_res1[12686],mul_res1[12687],mul_res1[12688],mul_res1[12689],mul_res1[12690],mul_res1[12691],mul_res1[12692],mul_res1[12693],mul_res1[12694],mul_res1[12695],mul_res1[12696],mul_res1[12697],mul_res1[12698],mul_res1[12699],mul_res1[12700],mul_res1[12701],mul_res1[12702],mul_res1[12703],mul_res1[12704],mul_res1[12705],mul_res1[12706],mul_res1[12707],mul_res1[12708],mul_res1[12709],mul_res1[12710],mul_res1[12711],mul_res1[12712],mul_res1[12713],mul_res1[12714],mul_res1[12715],mul_res1[12716],mul_res1[12717],mul_res1[12718],mul_res1[12719],mul_res1[12720],mul_res1[12721],mul_res1[12722],mul_res1[12723],mul_res1[12724],mul_res1[12725],mul_res1[12726],mul_res1[12727],mul_res1[12728],mul_res1[12729],mul_res1[12730],mul_res1[12731],mul_res1[12732],mul_res1[12733],mul_res1[12734],mul_res1[12735],mul_res1[12736],mul_res1[12737],mul_res1[12738],mul_res1[12739],mul_res1[12740],mul_res1[12741],mul_res1[12742],mul_res1[12743],mul_res1[12744],mul_res1[12745],mul_res1[12746],mul_res1[12747],mul_res1[12748],mul_res1[12749],mul_res1[12750],mul_res1[12751],mul_res1[12752],mul_res1[12753],mul_res1[12754],mul_res1[12755],mul_res1[12756],mul_res1[12757],mul_res1[12758],mul_res1[12759],mul_res1[12760],mul_res1[12761],mul_res1[12762],mul_res1[12763],mul_res1[12764],mul_res1[12765],mul_res1[12766],mul_res1[12767],mul_res1[12768],mul_res1[12769],mul_res1[12770],mul_res1[12771],mul_res1[12772],mul_res1[12773],mul_res1[12774],mul_res1[12775],mul_res1[12776],mul_res1[12777],mul_res1[12778],mul_res1[12779],mul_res1[12780],mul_res1[12781],mul_res1[12782],mul_res1[12783],mul_res1[12784],mul_res1[12785],mul_res1[12786],mul_res1[12787],mul_res1[12788],mul_res1[12789],mul_res1[12790],mul_res1[12791],mul_res1[12792],mul_res1[12793],mul_res1[12794],mul_res1[12795],mul_res1[12796],mul_res1[12797],mul_res1[12798],mul_res1[12799],result_fc1[63]);


  /*
  #include <stdio.h>  

void main() {
    int i = 0;
    int k=0;
    for (i = 0; i < 12800; i = i+200) {
        // Print the current element
        
        printf("adder_200in adder_200in_mod_%d(clk,rst,mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],mul_res1[%d],result_fc1[%d]);",k,i+0,i+1,i+2,i+3,i+4,i+5,i+6,i+7,i+8,i+9,i+10,i+11,i+12,i+13,i+14,i+15,i+16,i+17,i+18,i+19,i+20,i+21,i+22,i+23,i+24,i+25,i+26,i+27,i+28,i+29,i+30,i+31,i+32,i+33,i+34,i+35,i+36,i+37,i+38,i+39,i+40,i+41,i+42,i+43,i+44,i+45,i+46,i+47,i+48,i+49,i+50,i+51,i+52,i+53,i+54,i+55,i+56,i+57,i+58,i+59,i+60,i+61,i+62,i+63,i+64,i+65,i+66,i+67,i+68,i+69,i+70,i+71,i+72,i+73,i+74,i+75,i+76,i+77,i+78,i+79,i+80,i+81,i+82,i+83,i+84,i+85,i+86,i+87,i+88,i+89,i+90,i+91,i+92,i+93,i+94,i+95,i+96,i+97,i+98,i+99,i+100,i+101,i+102,i+103,i+104,i+105,i+106,i+107,i+108,i+109,i+110,i+111,i+112,i+113,i+114,i+115,i+116,i+117,i+118,i+119,i+120,i+121,i+122,i+123,i+124,i+125,i+126,i+127,i+128,i+129,i+130,i+131,i+132,i+133,i+134,i+135,i+136,i+137,i+138,i+139,i+140,i+141,i+142,i+143,i+144,i+145,i+146,i+147,i+148,i+149,i+150,i+151,i+152,i+153,i+154,i+155,i+156,i+157,i+158,i+159,i+160,i+161,i+162,i+163,i+164,i+165,i+166,i+167,i+168,i+169,i+170,i+171,i+172,i+173,i+174,i+175,i+176,i+177,i+178,i+179,i+180,i+181,i+182,i+183,i+184,i+185,i+186,i+187,i+188,i+189,i+190,i+191,i+192,i+193,i+194,i+195,i+196,i+197,i+198,i+199,k);  

        // Add a comma if it's not the last element in the current block of 200
       
            printf("\n\n\n");
            k = k+1;
        
    }
}
 
  
  
  
  
  */

integer k;
always_comb begin
        $write("matrix_B: ");
        foreach (matrix_B[k]) begin
            $write("%d, ", matrix_B[k]);  // Prints on the same line
        end
        $display("");  // Move to a new line after printing all values
    end


    
endmodule
